

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO square_root_finder 
  PIN rst 
    ANTENNAPARTIALMETALAREA 4.5626 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2727 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2232 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 23.453 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 90.8504 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.605735 LAYER VIA34 ;
  END rst
  PIN clk 
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.6432 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3032 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8529 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 20.4887 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 78.7263 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.237777 LAYER VIA45 ;
  END clk
  PIN in[15] 
    ANTENNAPARTIALMETALAREA 11.6788 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 44.2126 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.476 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0988 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 35.8904 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 136.464 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 121.478 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 466.171 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER VIA45 ;
  END in[15]
  PIN in[14] 
    ANTENNAPARTIALMETALAREA 13.2244 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 50.3606 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.724 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.6916 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 25.956 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 98.8556 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.54 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 52.0289 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 199.437 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 0.500741 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 5.2808 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.2884 LAYER METAL5 ;
    ANTENNAGATEAREA 0.648 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 60.1783 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 230.746 LAYER METAL5 ;
  END in[14]
  PIN in[13] 
    ANTENNAPARTIALMETALAREA 4.2252 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9954 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 8.0528 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.7824 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 39.676 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 150.499 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7344 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 64.3339 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 246.995 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.04321 LAYER VIA45 ;
  END in[13]
  PIN in[12] 
    ANTENNAPARTIALMETALAREA 16.6726 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.1177 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 32.9056 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 124.868 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 74.2929 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 283.485 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.834568 LAYER VIA45 ;
  END in[12]
  PIN in[11] 
    ANTENNAPARTIALMETALAREA 21.1526 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 80.0777 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 33.8744 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 128.536 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 62.3985 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 244.193 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER VIA45 ;
  END in[11]
  PIN in[10] 
    ANTENNAPARTIALMETALAREA 17.4552 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.0804 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 17.8304 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 68.0944 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 135.763 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 522.999 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 3.12963 LAYER VIA45 ;
  END in[10]
  PIN in[9] 
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 20.6682 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 79.4311 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0702 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 48.5732 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 186.915 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.17071 LAYER VIA45 ;
  END in[9]
  PIN in[8] 
    ANTENNAPARTIALMETALAREA 33.0806 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 125.531 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 64.2059 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 244.345 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.25185 LAYER VIA34 ;
  END in[8]
  PIN in[7] 
    ANTENNAPARTIALMETALAREA 47.152 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 179.098 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.54 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 90.3785 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 344.068 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.500741 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.2352 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1872 LAYER METAL4 ;
    ANTENNAGATEAREA 0.54 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 90.8141 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 346.267 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 0.625926 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 2.5088 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.7944 LAYER METAL5 ;
    ANTENNAGATEAREA 1.0702 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 93.1583 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 355.419 LAYER METAL5 ;
  END in[7]
  PIN in[6] 
    ANTENNAPARTIALMETALAREA 38.4636 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 145.612 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 11.1384 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 42.4636 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 24.325 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 97.9191 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER VIA45 ;
  END in[6]
  PIN in[5] 
    ANTENNAPARTIALMETALAREA 42.2086 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 159.79 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 20.2048 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 76.7864 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6696 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 51.4691 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 198.365 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.66577 LAYER VIA45 ;
  END in[5]
  PIN in[4] 
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.8276 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.787 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2232 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 37.0703 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 145.061 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.908602 LAYER VIA45 ;
  END in[4]
  PIN in[3] 
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2232 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 15.0067 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 67.746 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.605735 LAYER VIA34 ;
  END in[3]
  PIN in[2] 
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.5222 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2737 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2232 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 32.4225 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 127.466 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.908602 LAYER VIA45 ;
  END in[2]
  PIN in[1] 
    ANTENNAPARTIALMETALAREA 36.4406 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 137.954 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 54.8576 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 207.972 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 116.881 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 446.476 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.9821 LAYER VIA45 ;
  END in[1]
  PIN in[0] 
    ANTENNAPARTIALMETALAREA 38.9004 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 146.99 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 55.4848 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 210.346 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 1.1648 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5968 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 30.504 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 125.433 LAYER METAL5 ;
  END in[0]
  PIN sqrt[30] 
    ANTENNAPARTIALMETALAREA 2.75825 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.2131 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 38.7296 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 146.916 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 70.3836 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 267.639 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.2028 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 39.6816 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 151.114 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5972 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 40.6419 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 158.352 LAYER METAL5 ;
  END sqrt[30]
  PIN sqrt[29] 
    ANTENNAPARTIALMETALAREA 2.7272 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.3244 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 25.424 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 96.5448 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 75.5804 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 286.719 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.2704 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 48.2888 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 183.995 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7196 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 46.1255 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 177.837 LAYER METAL5 ;
  END sqrt[29]
  PIN sqrt[28] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.106 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.5532 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.7482 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.9568 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4904 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 53.256 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 204.283 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.112 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 137.722 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 529.926 LAYER METAL5 ;
  END sqrt[28]
  PIN sqrt[27] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.106 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.2078 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6549 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 74.3652 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 281.822 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 49.49 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 188.839 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2344 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 34.1332 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 130.104 LAYER METAL5 ;
  END sqrt[27]
  PIN sqrt[26] 
    ANTENNAPARTIALMETALAREA 0.028 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.106 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.2296 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.166 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 79.8252 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 302.492 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 33.74 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 128.027 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3568 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 91.0499 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 350.787 LAYER METAL5 ;
  END sqrt[26]
  PIN sqrt[25] 
    ANTENNAPARTIALMETALAREA 0.2772 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0494 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 29.4616 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 111.83 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 77.5852 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 294.012 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1268 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 112.278 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 429.391 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 1.24347 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 37.0664 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 140.62 LAYER METAL5 ;
    ANTENNAGATEAREA 2.7492 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 125.761 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 480.54 LAYER METAL5 ;
  END sqrt[25]
  PIN sqrt[24] 
    ANTENNAPARTIALMETALAREA 0.343 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2985 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 7.6832 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.3832 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 79.1308 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 300.457 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6224 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 81.4803 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 311.268 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 1.04315 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 40.9472 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 155.311 LAYER METAL5 ;
    ANTENNAGATEAREA 2.8716 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 123.674 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 474.818 LAYER METAL5 ;
  END sqrt[24]
  PIN sqrt[23] 
    ANTENNAPARTIALMETALAREA 0.3374 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2773 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.2072 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0812 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 86.1308 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 326.363 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 47.8128 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 181.896 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.994 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 147.733 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 565.386 LAYER METAL5 ;
  END sqrt[23]
  PIN sqrt[22] 
    ANTENNAPARTIALMETALAREA 1.8732 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0914 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 5.8352 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.3872 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.3888 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.5544 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 93.0384 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 353.998 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.1164 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 113.451 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 436.199 LAYER METAL5 ;
  END sqrt[22]
  PIN sqrt[21] 
    ANTENNAPARTIALMETALAREA 5.0302 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0429 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 62.0256 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 235.702 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8864 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 152.017 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 581.856 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.41067 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 28.14 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 106.827 LAYER METAL5 ;
    ANTENNAGATEAREA 3.7788 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 159.464 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 610.126 LAYER METAL5 ;
  END sqrt[21]
  PIN sqrt[20] 
    ANTENNAPARTIALMETALAREA 21.665 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 82.0175 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 52.9872 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 201.485 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0088 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 112.291 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 430.555 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 1.82859 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 15.8144 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 60.1656 LAYER METAL5 ;
    ANTENNAGATEAREA 3.9012 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 116.344 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 445.977 LAYER METAL5 ;
  END sqrt[20]
  PIN sqrt[19] 
    ANTENNAPARTIALMETALAREA 17.7856 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 67.3312 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 40.908 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 155.46 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0236 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 70.4936 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 273.959 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.71196 LAYER VIA45 ;
  END sqrt[19]
  PIN sqrt[18] 
    ANTENNAPARTIALMETALAREA 41.9258 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 160.203 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1016 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 138.712 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 530.067 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 1.71823 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 29.8032 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 113.42 LAYER METAL4 ;
    ANTENNAGATEAREA 4.146 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 145.9 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 557.424 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.72569 LAYER VIA45 ;
  END sqrt[18]
  PIN sqrt[17] 
    ANTENNADIFFAREA 1.2324 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 88.2546 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 337.075 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7284 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 86.1211 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 330.423 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 1.67499 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 21.7728 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 82.7224 LAYER METAL4 ;
    ANTENNAGATEAREA 4.2684 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 91.222 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 349.803 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.67499 LAYER VIA45 ;
  END sqrt[17]
  PIN sqrt[16] 
    ANTENNAPARTIALMETALAREA 7.9968 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.2736 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 47.04 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 179.564 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.3908 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 92.5279 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 355.431 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.27798 LAYER VIA45 ;
  END sqrt[16]
  PIN sqrt[15] 
    ANTENNAPARTIALMETALAREA 24.5756 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 93.333 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.54 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 78.7043 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 298.449 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.625926 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 70.6272 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 268.562 LAYER METAL4 ;
    ANTENNAGATEAREA 6.0108 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 134.895 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 516.131 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.29412 LAYER VIA45 ;
  END sqrt[15]
  PIN sqrt[14] 
    ANTENNAPARTIALMETALAREA 8.0206 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.3637 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNADIFFAREA 1.158 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 72.7356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 276.543 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.7832 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 72.7132 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 282.272 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.40738 LAYER VIA45 ;
    ANTENNADIFFAREA 1.158 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 20.2496 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 76.956 LAYER METAL5 ;
    ANTENNAGATEAREA 5.8632 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 76.1669 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 295.397 LAYER METAL5 ;
  END sqrt[14]
  PIN sqrt[13] 
    ANTENNAPARTIALMETALAREA 16.1504 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.1408 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 82.8912 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 315.286 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8232 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 134.442 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 522.74 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.30451 LAYER VIA45 ;
    ANTENNADIFFAREA 1.158 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 53.9896 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 204.983 LAYER METAL5 ;
    ANTENNAGATEAREA 5.9856 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 143.462 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 556.986 LAYER METAL5 ;
  END sqrt[13]
  PIN sqrt[12] 
    ANTENNAPARTIALMETALAREA 29.0836 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 110.102 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.2028 LAYER VIA34 ;
    ANTENNADIFFAREA 1.0164 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 104.236 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 396.684 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.1576 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 120.563 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 460.464 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.03816 LAYER VIA45 ;
    ANTENNADIFFAREA 1.0164 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 16.184 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 61.5648 LAYER METAL5 ;
    ANTENNAGATEAREA 6.2376 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 123.158 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 470.334 LAYER METAL5 ;
  END sqrt[12]
  PIN sqrt[11] 
    ANTENNAPARTIALMETALAREA 81.2238 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 308.084 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2096 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 73.336 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 278.941 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.487328 LAYER VIA34 ;
    ANTENNADIFFAREA 1.0164 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 80.9032 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 307.464 LAYER METAL4 ;
    ANTENNAGATEAREA 6.4896 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 121.674 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 465.176 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.84096 LAYER VIA45 ;
  END sqrt[11]
  PIN sqrt[10] 
    ANTENNAPARTIALMETALAREA 8.0122 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.3319 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 77.868 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 295.973 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.32 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 144.414 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 552.236 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.25844 LAYER VIA45 ;
  END sqrt[10]
  PIN sqrt[9] 
    ANTENNAPARTIALMETALAREA 3.0492 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4321 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 25.0432 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 95.4 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6696 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 47.3837 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 181.376 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 0.504779 LAYER VIA45 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 57.9488 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 219.674 LAYER METAL5 ;
    ANTENNAGATEAREA 7.0044 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 107.541 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 412.547 LAYER METAL5 ;
  END sqrt[9]
  PIN sqrt[8] 
    ANTENNAPARTIALMETALAREA 12.4278 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 47.3449 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 103.501 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 395.422 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA23 ;
    ANTENNAMAXCUTCAR 1.65686 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 79.8392 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 305.513 LAYER METAL3 ;
    ANTENNAGATEAREA 2.988 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 130.221 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 497.668 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.2704 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 1.74736 LAYER VIA34 ;
    ANTENNADIFFAREA 1.0164 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 63.1064 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 240.387 LAYER METAL4 ;
    ANTENNAGATEAREA 6.2412 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 140.332 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 536.184 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.20915 LAYER VIA45 ;
  END sqrt[8]
  PIN sqrt[7] 
    ANTENNAPARTIALMETALAREA 10.2004 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 38.6158 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 17.4776 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 66.462 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNADIFFAREA 3.9084 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 81.8496 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 311.343 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.18 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 86.3603 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 332.894 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.79493 LAYER VIA45 ;
  END sqrt[7]
  PIN sqrt[6] 
    ANTENNAPARTIALMETALAREA 13.6038 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 51.5001 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 63.7112 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 244.16 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3464 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 117.753 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 451.583 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.2028 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.35977 LAYER VIA34 ;
    ANTENNADIFFAREA 1.2324 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 42.0952 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 160.844 LAYER METAL4 ;
    ANTENNAGATEAREA 7.6308 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 123.27 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 472.661 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.35977 LAYER VIA45 ;
  END sqrt[6]
  PIN sqrt[5] 
    ANTENNAPARTIALMETALAREA 17.6792 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 67.2252 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 41.9272 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 160.802 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3464 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 93.5904 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 359.447 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.30957 LAYER VIA34 ;
    ANTENNADIFFAREA 2.321 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 39.48 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 150.647 LAYER METAL4 ;
    ANTENNAGATEAREA 7.4706 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 98.8751 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 379.612 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.30957 LAYER VIA45 ;
  END sqrt[5]
  PIN sqrt[4] 
    ANTENNAPARTIALMETALAREA 3.976 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.052 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNADIFFAREA 2.321 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 108.217 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 416.209 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.8048 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 115.489 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 442.165 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.23729 LAYER VIA34 ;
    ANTENNADIFFAREA 2.321 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 31.9256 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 122.048 LAYER METAL4 ;
    ANTENNAGATEAREA 8.826 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 119.106 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 455.994 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.23729 LAYER VIA45 ;
  END sqrt[4]
  PIN sqrt[3] 
    ANTENNAPARTIALMETALAREA 14.7126 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 55.6977 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA23 ;
    ANTENNADIFFAREA 6.5045 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 74.9056 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 287.43 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4584 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 81.8445 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 314.553 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.24824 LAYER VIA34 ;
    ANTENNADIFFAREA 6.5045 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 40.0736 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 152.598 LAYER METAL4 ;
    ANTENNAGATEAREA 9.4824 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 86.0706 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 330.645 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.24824 LAYER VIA45 ;
  END sqrt[3]
  PIN sqrt[2] 
    ANTENNAPARTIALMETALAREA 21.1288 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 79.9876 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.2028 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 40.236 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 154.4 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4688 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 56.8342 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 220.169 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 1.74891 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 10.276 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 39.4956 LAYER METAL4 ;
    ANTENNAGATEAREA 7.0764 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 85.6099 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 328.1 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 1.75846 LAYER VIA45 ;
    ANTENNADIFFAREA 6.5045 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 2.6936 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.494 LAYER METAL5 ;
    ANTENNAGATEAREA 9.678 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 85.8882 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 329.184 LAYER METAL5 ;
  END sqrt[2]
  PIN sqrt[1] 
    ANTENNAPARTIALMETALAREA 14.9422 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 56.5669 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNADIFFAREA 6.5045 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 38.5224 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 147.616 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6448 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 64.2249 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 254.997 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.23471 LAYER VIA34 ;
    ANTENNADIFFAREA 6.5045 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 8.5792 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.072 LAYER METAL4 ;
    ANTENNAGATEAREA 5.2152 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 89.4639 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 344.252 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.27471 LAYER VIA45 ;
    ANTENNADIFFAREA 6.5045 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 44.9064 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 170.596 LAYER METAL5 ;
    ANTENNAGATEAREA 10.4052 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 93.7796 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 360.647 LAYER METAL5 ;
  END sqrt[1]
  PIN sqrt[0] 
    ANTENNAPARTIALMETALAREA 3.6484 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8118 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA23 ;
    ANTENNADIFFAREA 5.2896 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 75.88 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 292.009 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.7944 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 101.929 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 398.119 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.24478 LAYER VIA34 ;
    ANTENNADIFFAREA 5.2896 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 38.598 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 146.715 LAYER METAL4 ;
    ANTENNAGATEAREA 9.8016 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 105.867 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 413.087 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.24478 LAYER VIA45 ;
  END sqrt[0]
END square_root_finder

END LIBRARY
