module square_root_finder();



endmodule
