
module square_root_finder_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;

  wire   [30:1] carry;

  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(SUM[31]), .S(
        SUM[30]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module square_root_finder_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;

  wire   [30:1] carry;

  ADDFX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFX2 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX2 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFX2 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFX2 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFX2 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  ADDFX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFX2 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  ADDFX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFX2 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFX2 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFX2 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFX2 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADDFX2 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFX2 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX2 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFX2 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX2 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFX2 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX2 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFX2 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX2 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFX2 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFX2 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFX2 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ADDFX2 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ADDFX2 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  ADDFX2 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(SUM[31]), .S(
        SUM[30]) );
  AND2X1 U1 ( .A(B[0]), .B(A[0]), .Y(carry[1]) );
endmodule


module square_root_finder_DW02_mult_2 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   ab_30__1_, ab_30__0_, ab_29__1_, ab_29__0_, ab_28__1_, ab_28__0_,
         ab_27__1_, ab_27__0_, ab_26__1_, ab_26__0_, ab_25__1_, ab_25__0_,
         ab_24__1_, ab_24__0_, ab_23__1_, ab_23__0_, ab_22__1_, ab_22__0_,
         ab_21__10_, ab_21__1_, ab_21__0_, ab_20__11_, ab_20__10_, ab_20__1_,
         ab_20__0_, ab_19__12_, ab_19__11_, ab_19__10_, ab_19__0_, ab_18__13_,
         ab_18__12_, ab_18__11_, ab_18__10_, ab_18__0_, ab_17__14_, ab_17__13_,
         ab_17__12_, ab_17__11_, ab_17__10_, ab_17__0_, ab_16__15_, ab_16__14_,
         ab_16__13_, ab_16__12_, ab_16__11_, ab_16__10_, ab_16__0_, ab_15__14_,
         ab_15__13_, ab_15__12_, ab_15__11_, ab_15__10_, ab_15__0_, ab_14__13_,
         ab_14__12_, ab_14__11_, ab_14__10_, ab_14__0_, ab_13__12_, ab_13__11_,
         ab_13__10_, ab_13__0_, ab_12__11_, ab_12__10_, ab_12__0_, ab_11__10_,
         ab_11__0_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_,
         ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_,
         ab_9__12_, ab_9__11_, ab_9__10_, ab_9__8_, ab_9__7_, ab_9__6_,
         ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__23_,
         ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_, ab_8__17_,
         ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_, ab_8__11_,
         ab_8__10_, ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_, ab_8__2_,
         ab_8__1_, ab_8__0_, ab_7__24_, ab_7__23_, ab_7__22_, ab_7__21_,
         ab_7__20_, ab_7__19_, ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_,
         ab_7__14_, ab_7__13_, ab_7__12_, ab_7__11_, ab_7__10_, ab_7__6_,
         ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__5_, ab_6__4_, ab_6__3_,
         ab_6__2_, ab_6__1_, ab_6__0_, ab_5__26_, ab_5__25_, ab_5__24_,
         ab_5__23_, ab_5__22_, ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_,
         ab_5__17_, ab_5__16_, ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_,
         ab_5__11_, ab_5__10_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_,
         ab_5__0_, ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_, ab_4__23_,
         ab_4__22_, ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_,
         ab_4__16_, ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_,
         ab_4__10_, ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__28_,
         ab_3__27_, ab_3__26_, ab_3__25_, ab_3__24_, ab_3__23_, ab_3__22_,
         ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_, ab_3__17_, ab_3__16_,
         ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_, ab_3__11_, ab_3__10_,
         ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_, ab_2__28_, ab_2__27_,
         ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_, ab_2__22_, ab_2__21_,
         ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_, ab_2__15_,
         ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_, ab_2__1_,
         ab_2__0_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_,
         ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, CARRYB_15__15_,
         CARRYB_15__14_, CARRYB_15__13_, CARRYB_15__12_, CARRYB_15__11_,
         CARRYB_15__10_, CARRYB_15__9_, CARRYB_15__8_, CARRYB_15__7_,
         CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_, CARRYB_15__3_,
         CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_, CARRYB_14__16_,
         CARRYB_14__15_, CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_,
         CARRYB_14__11_, CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_,
         CARRYB_14__7_, CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_,
         CARRYB_14__3_, CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_,
         CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_, CARRYB_13__14_,
         CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_, CARRYB_13__10_,
         CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_, CARRYB_13__6_,
         CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_,
         CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__18_, CARRYB_12__17_,
         CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_, CARRYB_12__13_,
         CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_, CARRYB_12__9_,
         CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_, CARRYB_12__5_,
         CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_,
         CARRYB_12__0_, CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_,
         CARRYB_11__16_, CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_,
         CARRYB_11__12_, CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_,
         CARRYB_11__8_, CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_,
         CARRYB_11__4_, CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_,
         CARRYB_11__0_, CARRYB_10__20_, CARRYB_10__19_, CARRYB_10__18_,
         CARRYB_10__17_, CARRYB_10__16_, CARRYB_10__15_, CARRYB_10__14_,
         CARRYB_10__13_, CARRYB_10__12_, CARRYB_10__11_, CARRYB_10__10_,
         CARRYB_10__9_, CARRYB_10__8_, CARRYB_10__7_, CARRYB_10__6_,
         CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_, CARRYB_10__2_,
         CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__21_, CARRYB_9__20_,
         CARRYB_9__19_, CARRYB_9__18_, CARRYB_9__17_, CARRYB_9__16_,
         CARRYB_9__15_, CARRYB_9__14_, CARRYB_9__13_, CARRYB_9__12_,
         CARRYB_9__11_, CARRYB_9__10_, CARRYB_9__9_, CARRYB_9__8_,
         CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_, CARRYB_9__4_, CARRYB_9__3_,
         CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_, CARRYB_8__22_,
         CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_, CARRYB_8__18_,
         CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_, CARRYB_8__14_,
         CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_, CARRYB_8__10_,
         CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_, CARRYB_8__5_,
         CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_, CARRYB_8__0_,
         CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_, CARRYB_7__20_,
         CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_, CARRYB_7__16_,
         CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_, CARRYB_7__12_,
         CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_, CARRYB_7__8_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, CARRYB_1__0_, SUMB_15__16_,
         SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_,
         SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_,
         SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_,
         SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_,
         SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_,
         SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_,
         SUMB_14__2_, SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__19_, SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_,
         SUMB_12__14_, SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_,
         SUMB_12__9_, SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_,
         SUMB_12__4_, SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_,
         SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_,
         SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_,
         SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_,
         SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_,
         SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_,
         SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_,
         SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_,
         SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_,
         SUMB_9__2_, SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__24_, SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_,
         SUMB_7__19_, SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_,
         SUMB_7__14_, SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_,
         SUMB_7__9_, SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_,
         SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_,
         SUMB_6__24_, SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_,
         SUMB_5__25_, SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_,
         SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_,
         SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_,
         SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_,
         SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_,
         SUMB_4__27_, SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_,
         SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_,
         SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_,
         SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_,
         SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_,
         SUMB_4__2_, SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_,
         SUMB_3__25_, SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__29_, SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_,
         SUMB_2__24_, SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_,
         SUMB_2__19_, SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_,
         SUMB_2__14_, SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_,
         SUMB_2__9_, SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_,
         SUMB_2__4_, SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__29_,
         SUMB_1__28_, SUMB_1__27_, SUMB_1__26_, SUMB_1__25_, SUMB_1__24_,
         SUMB_1__23_, SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_,
         SUMB_1__18_, SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_,
         SUMB_1__13_, SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_,
         SUMB_1__8_, SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_,
         SUMB_1__3_, SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_, CARRYB_29__1_,
         CARRYB_29__0_, CARRYB_28__2_, CARRYB_28__1_, CARRYB_28__0_,
         CARRYB_27__3_, CARRYB_27__2_, CARRYB_27__1_, CARRYB_27__0_,
         CARRYB_26__4_, CARRYB_26__3_, CARRYB_26__2_, CARRYB_26__1_,
         CARRYB_26__0_, CARRYB_25__5_, CARRYB_25__4_, CARRYB_25__3_,
         CARRYB_25__2_, CARRYB_25__1_, CARRYB_25__0_, CARRYB_24__6_,
         CARRYB_24__5_, CARRYB_24__4_, CARRYB_24__3_, CARRYB_24__2_,
         CARRYB_24__1_, CARRYB_24__0_, CARRYB_23__7_, CARRYB_23__6_,
         CARRYB_23__5_, CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_,
         CARRYB_23__1_, CARRYB_23__0_, CARRYB_22__8_, CARRYB_22__7_,
         CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_, CARRYB_22__3_,
         CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_, CARRYB_21__9_,
         CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_, CARRYB_21__5_,
         CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_, CARRYB_21__1_,
         CARRYB_21__0_, CARRYB_20__10_, CARRYB_20__9_, CARRYB_20__8_,
         CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_, CARRYB_20__4_,
         CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_, CARRYB_20__0_,
         CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_, CARRYB_19__8_,
         CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_, CARRYB_19__4_,
         CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_, CARRYB_19__0_,
         CARRYB_18__12_, CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_,
         CARRYB_18__8_, CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_,
         CARRYB_18__4_, CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_,
         CARRYB_18__0_, CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_,
         CARRYB_17__10_, CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_,
         CARRYB_17__6_, CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_,
         CARRYB_17__2_, CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__14_,
         CARRYB_16__13_, CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_,
         CARRYB_16__9_, CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_,
         CARRYB_16__5_, CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_,
         CARRYB_16__1_, CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_, SUMB_29__1_,
         SUMB_28__3_, SUMB_28__2_, SUMB_28__1_, SUMB_27__4_, SUMB_27__3_,
         SUMB_27__2_, SUMB_27__1_, SUMB_26__5_, SUMB_26__4_, SUMB_26__3_,
         SUMB_26__2_, SUMB_26__1_, SUMB_25__6_, SUMB_25__5_, SUMB_25__4_,
         SUMB_25__3_, SUMB_25__2_, SUMB_25__1_, SUMB_24__7_, SUMB_24__6_,
         SUMB_24__5_, SUMB_24__4_, SUMB_24__3_, SUMB_24__2_, SUMB_24__1_,
         SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_,
         SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_22__9_, SUMB_22__8_,
         SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_,
         SUMB_22__2_, SUMB_22__1_, SUMB_21__10_, SUMB_21__9_, SUMB_21__8_,
         SUMB_21__7_, SUMB_21__6_, SUMB_21__5_, SUMB_21__4_, SUMB_21__3_,
         SUMB_21__2_, SUMB_21__1_, SUMB_20__11_, SUMB_20__10_, SUMB_20__9_,
         SUMB_20__8_, SUMB_20__7_, SUMB_20__6_, SUMB_20__5_, SUMB_20__4_,
         SUMB_20__3_, SUMB_20__2_, SUMB_20__1_, SUMB_19__12_, SUMB_19__11_,
         SUMB_19__10_, SUMB_19__9_, SUMB_19__8_, SUMB_19__7_, SUMB_19__6_,
         SUMB_19__5_, SUMB_19__4_, SUMB_19__3_, SUMB_19__2_, SUMB_19__1_,
         SUMB_18__13_, SUMB_18__12_, SUMB_18__11_, SUMB_18__10_, SUMB_18__9_,
         SUMB_18__8_, SUMB_18__7_, SUMB_18__6_, SUMB_18__5_, SUMB_18__4_,
         SUMB_18__3_, SUMB_18__2_, SUMB_18__1_, SUMB_17__14_, SUMB_17__13_,
         SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_,
         SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_,
         SUMB_17__2_, SUMB_17__1_, SUMB_16__15_, SUMB_16__14_, SUMB_16__13_,
         SUMB_16__12_, SUMB_16__11_, SUMB_16__10_, SUMB_16__9_, SUMB_16__8_,
         SUMB_16__7_, SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_,
         SUMB_16__2_, SUMB_16__1_, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53;

  ADDFX2 S2_2_28 ( .A(ab_2__28_), .B(n32), .CI(SUMB_1__29_), .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  ADDFX2 S2_2_27 ( .A(ab_2__27_), .B(n31), .CI(SUMB_1__28_), .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  ADDFX2 S2_2_26 ( .A(ab_2__26_), .B(n30), .CI(SUMB_1__27_), .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  ADDFX2 S2_2_25 ( .A(ab_2__25_), .B(n29), .CI(SUMB_1__26_), .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  ADDFX2 S2_2_24 ( .A(ab_2__24_), .B(n28), .CI(SUMB_1__25_), .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  ADDFX2 S2_2_23 ( .A(ab_2__23_), .B(n27), .CI(SUMB_1__24_), .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  ADDFX2 S2_2_22 ( .A(ab_2__22_), .B(n26), .CI(SUMB_1__23_), .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  ADDFX2 S2_2_21 ( .A(ab_2__21_), .B(n25), .CI(SUMB_1__22_), .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  ADDFX2 S2_2_20 ( .A(ab_2__20_), .B(n24), .CI(SUMB_1__21_), .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  ADDFX2 S2_2_19 ( .A(ab_2__19_), .B(n23), .CI(SUMB_1__20_), .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  ADDFX2 S2_2_18 ( .A(ab_2__18_), .B(n22), .CI(SUMB_1__19_), .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  ADDFX2 S2_2_17 ( .A(ab_2__17_), .B(n21), .CI(SUMB_1__18_), .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  ADDFX2 S2_2_16 ( .A(ab_2__16_), .B(n20), .CI(SUMB_1__17_), .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  ADDFX2 S2_2_15 ( .A(ab_2__15_), .B(n19), .CI(SUMB_1__16_), .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  ADDFX2 S2_2_14 ( .A(ab_2__14_), .B(n18), .CI(SUMB_1__15_), .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  XOR3X2 S2_15_16 ( .A(ab_16__15_), .B(CARRYB_14__16_), .C(SUMB_14__17_), .Y(
        SUMB_15__16_) );
  XOR3X2 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .C(SUMB_15__16_), .Y(
        SUMB_16__15_) );
  XOR3X2 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .C(SUMB_16__15_), .Y(
        SUMB_17__14_) );
  XOR3X2 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .C(SUMB_17__14_), .Y(
        SUMB_18__13_) );
  XOR3X2 S2_11_20 ( .A(ab_20__11_), .B(CARRYB_10__20_), .C(SUMB_10__21_), .Y(
        SUMB_11__20_) );
  XOR3X2 S2_12_19 ( .A(ab_19__12_), .B(CARRYB_11__19_), .C(SUMB_11__20_), .Y(
        SUMB_12__19_) );
  XOR3X2 S2_13_18 ( .A(ab_18__13_), .B(CARRYB_12__18_), .C(SUMB_12__19_), .Y(
        SUMB_13__18_) );
  XOR3X2 S2_14_17 ( .A(ab_17__14_), .B(CARRYB_13__17_), .C(SUMB_13__18_), .Y(
        SUMB_14__17_) );
  XOR3X2 S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .C(SUMB_6__25_), .Y(
        SUMB_7__24_) );
  XOR3X2 S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .C(SUMB_7__24_), .Y(
        SUMB_8__23_) );
  XOR3X2 S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .C(SUMB_8__23_), .Y(
        SUMB_9__22_) );
  XOR3X2 S2_10_21 ( .A(ab_21__10_), .B(CARRYB_9__21_), .C(SUMB_9__22_), .Y(
        SUMB_10__21_) );
  XOR3X2 S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .C(SUMB_2__29_), .Y(
        SUMB_3__28_) );
  XOR3X2 S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .C(SUMB_3__28_), .Y(
        SUMB_4__27_) );
  XOR3X2 S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .C(SUMB_4__27_), .Y(
        SUMB_5__26_) );
  XOR3X2 S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .C(SUMB_5__26_), .Y(
        SUMB_6__25_) );
  XOR3X2 S2_2_29 ( .A(ab_2__29_), .B(n33), .C(ab_30__1_), .Y(SUMB_2__29_) );
  ADDFX2 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  ADDFX2 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  ADDFX2 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  ADDFX2 S2_14_16 ( .A(ab_16__14_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  ADDFX2 S2_13_17 ( .A(ab_17__13_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  ADDFX2 S2_13_16 ( .A(ab_16__13_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  ADDFX2 S2_12_18 ( .A(ab_18__12_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  ADDFX2 S2_12_17 ( .A(ab_17__12_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  ADDFX2 S2_12_16 ( .A(ab_16__12_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  ADDFX2 S2_11_19 ( .A(ab_19__11_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  ADDFX2 S2_11_18 ( .A(ab_18__11_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  ADDFX2 S2_11_17 ( .A(ab_17__11_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  ADDFX2 S2_11_16 ( .A(ab_16__11_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  ADDFX2 S2_10_20 ( .A(ab_20__10_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  ADDFX2 S2_10_19 ( .A(ab_19__10_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  ADDFX2 S2_10_18 ( .A(ab_18__10_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  ADDFX2 S2_10_17 ( .A(ab_17__10_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  ADDFX2 S2_10_16 ( .A(ab_16__10_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  ADDFX2 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  ADDFX2 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  ADDFX2 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  ADDFX2 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  ADDFX2 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  ADDFX2 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  ADDFX2 S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  ADDFX2 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  ADDFX2 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  ADDFX2 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  ADDFX2 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  ADDFX2 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  ADDFX2 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  ADDFX2 S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), .CO(
        CARRYB_7__23_), .S(SUMB_7__23_) );
  ADDFX2 S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  ADDFX2 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  ADDFX2 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  ADDFX2 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  ADDFX2 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  ADDFX2 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  ADDFX2 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  ADDFX2 S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), .CO(
        CARRYB_6__24_), .S(SUMB_6__24_) );
  ADDFX2 S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), .CO(
        CARRYB_6__23_), .S(SUMB_6__23_) );
  ADDFX2 S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  ADDFX2 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  ADDFX2 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  ADDFX2 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  ADDFX2 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  ADDFX2 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  ADDFX2 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  ADDFX2 S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), .CO(
        CARRYB_5__25_), .S(SUMB_5__25_) );
  ADDFX2 S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), .CO(
        CARRYB_5__24_), .S(SUMB_5__24_) );
  ADDFX2 S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), .CO(
        CARRYB_5__23_), .S(SUMB_5__23_) );
  ADDFX2 S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  ADDFX2 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  ADDFX2 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  ADDFX2 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  ADDFX2 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  ADDFX2 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  ADDFX2 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  ADDFX2 S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), .CO(
        CARRYB_4__26_), .S(SUMB_4__26_) );
  ADDFX2 S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), .CO(
        CARRYB_4__25_), .S(SUMB_4__25_) );
  ADDFX2 S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), .CO(
        CARRYB_4__24_), .S(SUMB_4__24_) );
  ADDFX2 S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), .CO(
        CARRYB_4__23_), .S(SUMB_4__23_) );
  ADDFX2 S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  ADDFX2 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  ADDFX2 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  ADDFX2 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  ADDFX2 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  ADDFX2 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  ADDFX2 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  ADDFX2 S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), .CO(
        CARRYB_3__27_), .S(SUMB_3__27_) );
  ADDFX2 S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), .CO(
        CARRYB_3__26_), .S(SUMB_3__26_) );
  ADDFX2 S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), .CO(
        CARRYB_3__25_), .S(SUMB_3__25_) );
  ADDFX2 S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), .CO(
        CARRYB_3__24_), .S(SUMB_3__24_) );
  ADDFX2 S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), .CO(
        CARRYB_3__23_), .S(SUMB_3__23_) );
  ADDFX2 S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  ADDFX2 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  ADDFX2 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  ADDFX2 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  ADDFX2 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  ADDFX2 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  ADDFX2 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  ADDFX2 S2_15_15 ( .A(B[15]), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  ADDFX2 S2_14_14 ( .A(B[14]), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  ADDFX2 S2_13_13 ( .A(B[13]), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  XOR3X2 S2_23_8 ( .A(ab_8__23_), .B(CARRYB_22__8_), .C(SUMB_22__9_), .Y(
        SUMB_23__8_) );
  XOR3X2 S2_24_7 ( .A(ab_7__24_), .B(CARRYB_23__7_), .C(SUMB_23__8_), .Y(
        SUMB_24__7_) );
  XOR3X2 S2_25_6 ( .A(ab_6__25_), .B(CARRYB_24__6_), .C(SUMB_24__7_), .Y(
        SUMB_25__6_) );
  XOR3X2 S2_26_5 ( .A(ab_5__26_), .B(CARRYB_25__5_), .C(SUMB_25__6_), .Y(
        SUMB_26__5_) );
  XOR3X2 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .C(SUMB_18__13_), .Y(
        SUMB_19__12_) );
  XOR3X2 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .C(SUMB_19__12_), .Y(
        SUMB_20__11_) );
  XOR3X2 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .C(SUMB_20__11_), .Y(
        SUMB_21__10_) );
  XOR3X2 S2_22_9 ( .A(ab_9__22_), .B(CARRYB_21__9_), .C(SUMB_21__10_), .Y(
        SUMB_22__9_) );
  ADDFX2 S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), .CO(
        CARRYB_30__0_), .S(PRODUCT[30]) );
  ADDFX2 S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), .CO(
        CARRYB_27__0_), .S(PRODUCT[27]) );
  ADDFX2 S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), .CO(
        CARRYB_28__0_), .S(PRODUCT[28]) );
  ADDFX2 S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), .CO(
        CARRYB_29__0_), .S(PRODUCT[29]) );
  ADDFX2 S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), .CO(
        CARRYB_26__0_), .S(PRODUCT[26]) );
  ADDFX2 S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), .CO(
        CARRYB_25__0_), .S(PRODUCT[25]) );
  ADDFX2 S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), .CO(
        CARRYB_24__0_), .S(PRODUCT[24]) );
  ADDFX2 S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(PRODUCT[23]) );
  ADDFX2 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(PRODUCT[22]) );
  ADDFX2 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(PRODUCT[21]) );
  ADDFX2 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(PRODUCT[20]) );
  ADDFX2 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(PRODUCT[19]) );
  ADDFX2 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(PRODUCT[18]) );
  ADDFX2 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(PRODUCT[17]) );
  ADDFX2 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(PRODUCT[16]) );
  ADDFX2 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(SUMB_1__1_), .CO(
        CARRYB_2__0_), .S() );
  ADDFX2 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S() );
  ADDFX2 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S() );
  ADDFX2 S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), .CO(
        CARRYB_29__1_), .S(SUMB_29__1_) );
  ADDFX2 S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), .CO(
        CARRYB_28__1_), .S(SUMB_28__1_) );
  ADDFX2 S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), .CO(
        CARRYB_27__1_), .S(SUMB_27__1_) );
  ADDFX2 S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), .CO(
        CARRYB_26__1_), .S(SUMB_26__1_) );
  ADDFX2 S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), .CO(
        CARRYB_25__1_), .S(SUMB_25__1_) );
  ADDFX2 S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), .CO(
        CARRYB_24__1_), .S(SUMB_24__1_) );
  ADDFX2 S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  ADDFX2 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  ADDFX2 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  ADDFX2 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  ADDFX2 S2_19_1 ( .A(ab_1__19_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  ADDFX2 S2_18_1 ( .A(ab_1__18_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  ADDFX2 S2_17_1 ( .A(ab_1__17_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  ADDFX2 S2_16_1 ( .A(ab_1__16_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFX2 S2_28_2 ( .A(ab_2__28_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), .CO(
        CARRYB_28__2_), .S(SUMB_28__2_) );
  ADDFX2 S2_27_3 ( .A(ab_3__27_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), .CO(
        CARRYB_27__3_), .S(SUMB_27__3_) );
  ADDFX2 S2_27_2 ( .A(ab_2__27_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), .CO(
        CARRYB_27__2_), .S(SUMB_27__2_) );
  ADDFX2 S2_26_4 ( .A(ab_4__26_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), .CO(
        CARRYB_26__4_), .S(SUMB_26__4_) );
  ADDFX2 S2_26_3 ( .A(ab_3__26_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), .CO(
        CARRYB_26__3_), .S(SUMB_26__3_) );
  ADDFX2 S2_26_2 ( .A(ab_2__26_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), .CO(
        CARRYB_26__2_), .S(SUMB_26__2_) );
  ADDFX2 S2_25_5 ( .A(ab_5__25_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), .CO(
        CARRYB_25__5_), .S(SUMB_25__5_) );
  ADDFX2 S2_25_4 ( .A(ab_4__25_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), .CO(
        CARRYB_25__4_), .S(SUMB_25__4_) );
  ADDFX2 S2_25_3 ( .A(ab_3__25_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), .CO(
        CARRYB_25__3_), .S(SUMB_25__3_) );
  ADDFX2 S2_25_2 ( .A(ab_2__25_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), .CO(
        CARRYB_25__2_), .S(SUMB_25__2_) );
  ADDFX2 S2_24_6 ( .A(ab_6__24_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), .CO(
        CARRYB_24__6_), .S(SUMB_24__6_) );
  ADDFX2 S2_24_5 ( .A(ab_5__24_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), .CO(
        CARRYB_24__5_), .S(SUMB_24__5_) );
  ADDFX2 S2_24_4 ( .A(ab_4__24_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), .CO(
        CARRYB_24__4_), .S(SUMB_24__4_) );
  ADDFX2 S2_24_3 ( .A(ab_3__24_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), .CO(
        CARRYB_24__3_), .S(SUMB_24__3_) );
  ADDFX2 S2_24_2 ( .A(ab_2__24_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), .CO(
        CARRYB_24__2_), .S(SUMB_24__2_) );
  ADDFX2 S2_23_7 ( .A(ab_7__23_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  ADDFX2 S2_23_6 ( .A(ab_6__23_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  ADDFX2 S2_23_5 ( .A(ab_5__23_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  ADDFX2 S2_23_4 ( .A(ab_4__23_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  ADDFX2 S2_23_3 ( .A(ab_3__23_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  ADDFX2 S2_23_2 ( .A(ab_2__23_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  ADDFX2 S2_22_8 ( .A(ab_8__22_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  ADDFX2 S2_22_7 ( .A(ab_7__22_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  ADDFX2 S2_22_6 ( .A(ab_6__22_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  ADDFX2 S2_22_5 ( .A(ab_5__22_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  ADDFX2 S2_22_4 ( .A(ab_4__22_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  ADDFX2 S2_22_3 ( .A(ab_3__22_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  ADDFX2 S2_22_2 ( .A(ab_2__22_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  ADDFX2 S2_21_9 ( .A(ab_9__21_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  ADDFX2 S2_21_8 ( .A(ab_8__21_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  ADDFX2 S2_21_7 ( .A(ab_7__21_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  ADDFX2 S2_21_6 ( .A(ab_6__21_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  ADDFX2 S2_21_5 ( .A(ab_5__21_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  ADDFX2 S2_21_4 ( .A(ab_4__21_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  ADDFX2 S2_21_3 ( .A(ab_3__21_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  ADDFX2 S2_21_2 ( .A(ab_2__21_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  ADDFX2 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  ADDFX2 S2_20_9 ( .A(ab_9__20_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  ADDFX2 S2_20_8 ( .A(ab_8__20_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  ADDFX2 S2_20_7 ( .A(ab_7__20_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  ADDFX2 S2_20_6 ( .A(ab_6__20_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  ADDFX2 S2_20_5 ( .A(ab_5__20_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  ADDFX2 S2_20_4 ( .A(ab_4__20_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  ADDFX2 S2_20_3 ( .A(ab_3__20_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  ADDFX2 S2_20_2 ( .A(ab_2__20_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  ADDFX2 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  ADDFX2 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  ADDFX2 S2_19_9 ( .A(ab_9__19_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  ADDFX2 S2_19_8 ( .A(ab_8__19_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  ADDFX2 S2_19_7 ( .A(ab_7__19_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  ADDFX2 S2_19_6 ( .A(ab_6__19_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  ADDFX2 S2_19_5 ( .A(ab_5__19_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  ADDFX2 S2_19_4 ( .A(ab_4__19_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  ADDFX2 S2_19_3 ( .A(ab_3__19_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  ADDFX2 S2_19_2 ( .A(ab_2__19_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  ADDFX2 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  ADDFX2 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  ADDFX2 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  ADDFX2 S2_18_9 ( .A(ab_9__18_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  ADDFX2 S2_18_8 ( .A(ab_8__18_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  ADDFX2 S2_18_7 ( .A(ab_7__18_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  ADDFX2 S2_18_6 ( .A(ab_6__18_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  ADDFX2 S2_18_5 ( .A(ab_5__18_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  ADDFX2 S2_18_4 ( .A(ab_4__18_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  ADDFX2 S2_18_3 ( .A(ab_3__18_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  ADDFX2 S2_18_2 ( .A(ab_2__18_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  ADDFX2 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  ADDFX2 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  ADDFX2 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  ADDFX2 S2_17_9 ( .A(ab_9__17_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  ADDFX2 S2_17_8 ( .A(ab_8__17_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  ADDFX2 S2_17_7 ( .A(ab_7__17_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  ADDFX2 S2_17_6 ( .A(ab_6__17_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  ADDFX2 S2_17_5 ( .A(ab_5__17_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  ADDFX2 S2_17_4 ( .A(ab_4__17_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  ADDFX2 S2_17_3 ( .A(ab_3__17_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  ADDFX2 S2_17_2 ( .A(ab_2__17_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  ADDFX2 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  ADDFX2 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  ADDFX2 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  ADDFX2 S2_16_9 ( .A(ab_9__16_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  ADDFX2 S2_16_8 ( .A(ab_8__16_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  ADDFX2 S2_16_7 ( .A(ab_7__16_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  ADDFX2 S2_16_6 ( .A(ab_6__16_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFX2 S2_16_5 ( .A(ab_5__16_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFX2 S2_16_4 ( .A(ab_4__16_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFX2 S2_16_3 ( .A(ab_3__16_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFX2 S2_16_2 ( .A(ab_2__16_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  XOR3X2 S2_27_4 ( .A(ab_4__27_), .B(CARRYB_26__4_), .C(SUMB_26__5_), .Y(
        SUMB_27__4_) );
  XOR3X2 S2_28_3 ( .A(ab_3__28_), .B(CARRYB_27__3_), .C(SUMB_27__4_), .Y(
        SUMB_28__3_) );
  XOR3X2 S2_29_2 ( .A(ab_2__29_), .B(CARRYB_28__2_), .C(SUMB_28__3_), .Y(
        SUMB_29__2_) );
  XOR3X2 S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .C(SUMB_29__2_), .Y(
        SUMB_30__1_) );
  ADDFX2 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  ADDFX2 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  ADDFX2 S2_14_15 ( .A(ab_15__14_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  ADDFX2 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  ADDFX2 S2_13_15 ( .A(ab_15__13_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  ADDFX2 S2_13_14 ( .A(ab_14__13_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  ADDFX2 S2_12_15 ( .A(ab_15__12_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  ADDFX2 S2_12_14 ( .A(ab_14__12_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  ADDFX2 S2_12_13 ( .A(ab_13__12_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  ADDFX2 S2_11_15 ( .A(ab_15__11_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  ADDFX2 S2_11_14 ( .A(ab_14__11_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  ADDFX2 S2_11_13 ( .A(ab_13__11_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  ADDFX2 S2_10_15 ( .A(ab_15__10_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  ADDFX2 S2_10_14 ( .A(ab_14__10_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  ADDFX2 S2_10_13 ( .A(ab_13__10_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  ADDFX2 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  ADDFX2 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  ADDFX2 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  ADDFX2 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  ADDFX2 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  ADDFX2 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  ADDFX2 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  ADDFX2 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  ADDFX2 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  ADDFX2 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  ADDFX2 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  ADDFX2 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  ADDFX2 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  ADDFX2 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  ADDFX2 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  ADDFX2 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  ADDFX2 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  ADDFX2 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  ADDFX2 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  ADDFX2 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  ADDFX2 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  ADDFX2 S2_2_9 ( .A(ab_9__2_), .B(n15), .CI(SUMB_1__10_), .CO(CARRYB_2__9_), 
        .S(SUMB_2__9_) );
  ADDFX2 S2_2_8 ( .A(ab_8__2_), .B(n14), .CI(SUMB_1__9_), .CO(CARRYB_2__8_), 
        .S(SUMB_2__8_) );
  ADDFX2 S2_2_4 ( .A(ab_4__2_), .B(n10), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFX2 S2_2_3 ( .A(ab_3__2_), .B(n9), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFX2 S2_2_13 ( .A(ab_2__13_), .B(n17), .CI(SUMB_1__14_), .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  ADDFX2 S2_2_12 ( .A(ab_2__12_), .B(n16), .CI(SUMB_1__13_), .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  ADDFX2 S2_2_11 ( .A(ab_2__11_), .B(n13), .CI(SUMB_1__12_), .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  ADDFX2 S2_2_10 ( .A(ab_2__10_), .B(n12), .CI(SUMB_1__11_), .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  ADDFX2 S2_2_7 ( .A(ab_7__2_), .B(n11), .CI(SUMB_1__8_), .CO(CARRYB_2__7_), 
        .S(SUMB_2__7_) );
  ADDFX2 S2_2_6 ( .A(ab_6__2_), .B(n8), .CI(SUMB_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFX2 S2_2_5 ( .A(ab_5__2_), .B(n7), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFX2 S2_2_2 ( .A(n36), .B(n6), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  ADDFX2 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(PRODUCT[15]) );
  ADDFX2 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(PRODUCT[14]) );
  ADDFX2 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(PRODUCT[13]) );
  ADDFX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S() );
  ADDFX2 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S() );
  ADDFX2 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S() );
  ADDFX2 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(PRODUCT[12]) );
  ADDFX2 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S() );
  ADDFX2 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S() );
  ADDFX2 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S() );
  ADDFX2 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S() );
  ADDFX2 S2_15_1 ( .A(ab_1__15_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFX2 S2_14_1 ( .A(ab_1__14_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFX2 S2_13_1 ( .A(ab_1__13_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFX2 S2_2_1 ( .A(ab_2__1_), .B(n5), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFX2 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  ADDFX2 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  ADDFX2 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  ADDFX2 S2_15_9 ( .A(ab_9__15_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  ADDFX2 S2_15_8 ( .A(ab_8__15_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  ADDFX2 S2_15_7 ( .A(ab_7__15_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  ADDFX2 S2_15_6 ( .A(ab_6__15_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFX2 S2_15_5 ( .A(ab_5__15_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFX2 S2_15_4 ( .A(ab_4__15_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFX2 S2_15_3 ( .A(ab_3__15_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFX2 S2_15_2 ( .A(ab_2__15_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFX2 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  ADDFX2 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  ADDFX2 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  ADDFX2 S2_14_9 ( .A(ab_9__14_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  ADDFX2 S2_14_8 ( .A(ab_8__14_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  ADDFX2 S2_14_7 ( .A(ab_7__14_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  ADDFX2 S2_14_6 ( .A(ab_6__14_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFX2 S2_14_5 ( .A(ab_5__14_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFX2 S2_14_4 ( .A(ab_4__14_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFX2 S2_14_3 ( .A(ab_3__14_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFX2 S2_14_2 ( .A(ab_2__14_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFX2 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  ADDFX2 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  ADDFX2 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  ADDFX2 S2_13_9 ( .A(ab_9__13_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  ADDFX2 S2_13_8 ( .A(ab_8__13_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  ADDFX2 S2_13_7 ( .A(ab_7__13_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  ADDFX2 S2_13_6 ( .A(ab_6__13_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFX2 S2_13_5 ( .A(ab_5__13_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFX2 S2_13_4 ( .A(ab_4__13_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFX2 S2_13_3 ( .A(ab_3__13_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFX2 S2_13_2 ( .A(ab_2__13_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFX2 S2_12_12 ( .A(A[12]), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  ADDFX2 S2_11_11 ( .A(n52), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  ADDFX2 S2_10_10 ( .A(n50), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  ADDFX2 S2_9_9 ( .A(A[9]), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  ADDFX2 S2_8_8 ( .A(n48), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(CARRYB_8__8_), .S(SUMB_8__8_) );
  ADDFX2 S2_7_7 ( .A(n46), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(CARRYB_7__7_), .S(SUMB_7__7_) );
  ADDFX2 S2_6_6 ( .A(n44), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFX2 S2_5_5 ( .A(n42), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFX2 S2_4_4 ( .A(n40), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFX2 S2_3_3 ( .A(n38), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFX2 S2_12_1 ( .A(ab_1__12_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFX2 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFX2 S2_11_1 ( .A(ab_1__11_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFX2 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFX2 S2_10_1 ( .A(ab_1__10_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFX2 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFX2 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFX2 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFX2 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFX2 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  ADDFX2 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  ADDFX2 S2_12_9 ( .A(ab_9__12_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  ADDFX2 S2_12_8 ( .A(ab_8__12_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  ADDFX2 S2_12_7 ( .A(ab_7__12_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  ADDFX2 S2_12_6 ( .A(ab_6__12_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFX2 S2_12_5 ( .A(ab_5__12_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFX2 S2_12_4 ( .A(ab_4__12_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFX2 S2_12_3 ( .A(ab_3__12_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFX2 S2_12_2 ( .A(ab_2__12_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFX2 S2_11_12 ( .A(ab_12__11_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  ADDFX2 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  ADDFX2 S2_11_9 ( .A(ab_9__11_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  ADDFX2 S2_11_8 ( .A(ab_8__11_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  ADDFX2 S2_11_7 ( .A(ab_7__11_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  ADDFX2 S2_11_6 ( .A(ab_6__11_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFX2 S2_11_5 ( .A(ab_5__11_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFX2 S2_11_4 ( .A(ab_4__11_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFX2 S2_11_3 ( .A(ab_3__11_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFX2 S2_11_2 ( .A(ab_2__11_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFX2 S2_10_12 ( .A(ab_12__10_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  ADDFX2 S2_10_11 ( .A(ab_11__10_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  ADDFX2 S2_10_9 ( .A(ab_9__10_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  ADDFX2 S2_10_8 ( .A(ab_8__10_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  ADDFX2 S2_10_7 ( .A(ab_7__10_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  ADDFX2 S2_10_6 ( .A(ab_6__10_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFX2 S2_10_5 ( .A(ab_5__10_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFX2 S2_10_4 ( .A(ab_4__10_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFX2 S2_10_3 ( .A(ab_3__10_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFX2 S2_10_2 ( .A(ab_2__10_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFX2 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  ADDFX2 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  ADDFX2 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  ADDFX2 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  ADDFX2 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  ADDFX2 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFX2 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFX2 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFX2 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFX2 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFX2 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  ADDFX2 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  ADDFX2 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  ADDFX2 S2_8_9 ( .A(ab_9__8_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  ADDFX2 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  ADDFX2 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFX2 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFX2 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFX2 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFX2 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  ADDFX2 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  ADDFX2 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  ADDFX2 S2_7_9 ( .A(ab_9__7_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  ADDFX2 S2_7_8 ( .A(ab_8__7_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  ADDFX2 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFX2 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFX2 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFX2 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFX2 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFX2 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  ADDFX2 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  ADDFX2 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  ADDFX2 S2_6_9 ( .A(ab_9__6_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  ADDFX2 S2_6_8 ( .A(ab_8__6_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  ADDFX2 S2_6_7 ( .A(ab_7__6_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  ADDFX2 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFX2 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFX2 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFX2 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFX2 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  ADDFX2 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  ADDFX2 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  ADDFX2 S2_5_9 ( .A(ab_9__5_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  ADDFX2 S2_5_8 ( .A(ab_8__5_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  ADDFX2 S2_5_7 ( .A(ab_7__5_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  ADDFX2 S2_5_6 ( .A(ab_6__5_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFX2 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFX2 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  ADDFX2 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  ADDFX2 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  ADDFX2 S2_4_9 ( .A(ab_9__4_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  ADDFX2 S2_4_8 ( .A(ab_8__4_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  ADDFX2 S2_4_7 ( .A(ab_7__4_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  ADDFX2 S2_4_6 ( .A(ab_6__4_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFX2 S2_4_5 ( .A(ab_5__4_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFX2 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFX2 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFX2 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  ADDFX2 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  ADDFX2 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  ADDFX2 S2_3_9 ( .A(ab_9__3_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  ADDFX2 S2_3_8 ( .A(ab_8__3_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  ADDFX2 S2_3_7 ( .A(ab_7__3_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  ADDFX2 S2_3_6 ( .A(ab_6__3_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFX2 S2_3_5 ( .A(ab_5__3_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFX2 S2_3_4 ( .A(ab_4__3_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFX2 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  AND2X2 U2 ( .A(ab_2__0_), .B(n34), .Y(n5) );
  AND2X2 U3 ( .A(ab_3__0_), .B(ab_2__1_), .Y(n6) );
  AND2X2 U4 ( .A(ab_6__0_), .B(ab_5__1_), .Y(n7) );
  AND2X2 U5 ( .A(ab_7__0_), .B(ab_6__1_), .Y(n8) );
  AND2X2 U6 ( .A(ab_4__0_), .B(ab_3__1_), .Y(n9) );
  AND2X2 U7 ( .A(ab_5__0_), .B(ab_4__1_), .Y(n10) );
  AND2X2 U8 ( .A(ab_8__0_), .B(ab_7__1_), .Y(n11) );
  AND2X2 U9 ( .A(ab_11__0_), .B(ab_1__10_), .Y(n12) );
  AND2X2 U10 ( .A(ab_12__0_), .B(ab_1__11_), .Y(n13) );
  AND2X2 U11 ( .A(ab_9__0_), .B(ab_8__1_), .Y(n14) );
  AND2X2 U12 ( .A(ab_10__0_), .B(ab_9__1_), .Y(n15) );
  AND2X2 U13 ( .A(ab_13__0_), .B(ab_1__12_), .Y(n16) );
  AND2X2 U14 ( .A(ab_14__0_), .B(ab_1__13_), .Y(n17) );
  AND2X2 U15 ( .A(ab_15__0_), .B(ab_1__14_), .Y(n18) );
  AND2X2 U16 ( .A(ab_16__0_), .B(ab_1__15_), .Y(n19) );
  AND2X2 U17 ( .A(ab_17__0_), .B(ab_1__16_), .Y(n20) );
  AND2X2 U18 ( .A(ab_18__0_), .B(ab_1__17_), .Y(n21) );
  AND2X2 U19 ( .A(ab_19__0_), .B(ab_1__18_), .Y(n22) );
  AND2X2 U20 ( .A(ab_20__0_), .B(ab_1__19_), .Y(n23) );
  AND2X2 U21 ( .A(ab_21__0_), .B(ab_20__1_), .Y(n24) );
  AND2X2 U22 ( .A(ab_22__0_), .B(ab_21__1_), .Y(n25) );
  AND2X2 U23 ( .A(ab_23__0_), .B(ab_22__1_), .Y(n26) );
  AND2X2 U24 ( .A(ab_24__0_), .B(ab_23__1_), .Y(n27) );
  AND2X2 U25 ( .A(ab_25__0_), .B(ab_24__1_), .Y(n28) );
  AND2X2 U26 ( .A(ab_26__0_), .B(ab_25__1_), .Y(n29) );
  AND2X2 U27 ( .A(ab_27__0_), .B(ab_26__1_), .Y(n30) );
  AND2X2 U28 ( .A(ab_28__0_), .B(ab_27__1_), .Y(n31) );
  AND2X2 U29 ( .A(ab_29__0_), .B(ab_28__1_), .Y(n32) );
  AND2X2 U30 ( .A(ab_30__0_), .B(ab_29__1_), .Y(n33) );
  XOR2X1 U31 ( .A(ab_2__1_), .B(ab_3__0_), .Y(SUMB_1__2_) );
  XOR2X1 U32 ( .A(ab_3__1_), .B(ab_4__0_), .Y(SUMB_1__3_) );
  XOR2X1 U33 ( .A(ab_6__1_), .B(ab_7__0_), .Y(SUMB_1__6_) );
  XOR2X1 U34 ( .A(ab_7__1_), .B(ab_8__0_), .Y(SUMB_1__7_) );
  XOR2X1 U35 ( .A(ab_8__1_), .B(ab_9__0_), .Y(SUMB_1__8_) );
  XOR2X1 U36 ( .A(ab_1__11_), .B(ab_12__0_), .Y(SUMB_1__11_) );
  XOR2X1 U37 ( .A(ab_1__12_), .B(ab_13__0_), .Y(SUMB_1__12_) );
  XOR2X1 U38 ( .A(ab_1__13_), .B(ab_14__0_), .Y(SUMB_1__13_) );
  XOR2X1 U39 ( .A(ab_1__14_), .B(ab_15__0_), .Y(SUMB_1__14_) );
  XOR2X1 U40 ( .A(ab_4__1_), .B(ab_5__0_), .Y(SUMB_1__4_) );
  XOR2X1 U41 ( .A(ab_5__1_), .B(ab_6__0_), .Y(SUMB_1__5_) );
  XOR2X1 U42 ( .A(ab_9__1_), .B(ab_10__0_), .Y(SUMB_1__9_) );
  XOR2X1 U43 ( .A(ab_1__10_), .B(ab_11__0_), .Y(SUMB_1__10_) );
  XOR2X1 U44 ( .A(n34), .B(ab_2__0_), .Y(SUMB_1__1_) );
  INVX1 U45 ( .A(n41), .Y(n40) );
  INVX1 U46 ( .A(B[4]), .Y(n41) );
  INVX1 U47 ( .A(n43), .Y(n42) );
  INVX1 U48 ( .A(B[5]), .Y(n43) );
  INVX1 U49 ( .A(n45), .Y(n44) );
  INVX1 U50 ( .A(B[6]), .Y(n45) );
  INVX1 U51 ( .A(n47), .Y(n46) );
  INVX1 U52 ( .A(B[7]), .Y(n47) );
  INVX1 U53 ( .A(n49), .Y(n48) );
  INVX1 U54 ( .A(B[8]), .Y(n49) );
  INVX1 U55 ( .A(n37), .Y(n36) );
  INVX1 U56 ( .A(B[2]), .Y(n37) );
  INVX1 U57 ( .A(n39), .Y(n38) );
  INVX1 U58 ( .A(B[3]), .Y(n39) );
  INVX1 U59 ( .A(n35), .Y(n34) );
  INVX1 U60 ( .A(B[1]), .Y(n35) );
  INVX1 U61 ( .A(n51), .Y(n50) );
  INVX1 U62 ( .A(B[10]), .Y(n51) );
  INVX1 U63 ( .A(n53), .Y(n52) );
  INVX1 U64 ( .A(B[11]), .Y(n53) );
  XOR2X1 U65 ( .A(ab_1__15_), .B(ab_16__0_), .Y(SUMB_1__15_) );
  XOR2X1 U66 ( .A(ab_1__16_), .B(ab_17__0_), .Y(SUMB_1__16_) );
  XOR2X1 U67 ( .A(ab_1__17_), .B(ab_18__0_), .Y(SUMB_1__17_) );
  XOR2X1 U68 ( .A(ab_1__18_), .B(ab_19__0_), .Y(SUMB_1__18_) );
  XOR2X1 U69 ( .A(ab_1__19_), .B(ab_20__0_), .Y(SUMB_1__19_) );
  XOR2X1 U70 ( .A(ab_20__1_), .B(ab_21__0_), .Y(SUMB_1__20_) );
  XOR2X1 U71 ( .A(ab_21__1_), .B(ab_22__0_), .Y(SUMB_1__21_) );
  XOR2X1 U72 ( .A(ab_22__1_), .B(ab_23__0_), .Y(SUMB_1__22_) );
  XOR2X1 U73 ( .A(ab_23__1_), .B(ab_24__0_), .Y(SUMB_1__23_) );
  XOR2X1 U74 ( .A(ab_24__1_), .B(ab_25__0_), .Y(SUMB_1__24_) );
  XOR2X1 U75 ( .A(ab_25__1_), .B(ab_26__0_), .Y(SUMB_1__25_) );
  XOR2X1 U76 ( .A(ab_26__1_), .B(ab_27__0_), .Y(SUMB_1__26_) );
  XOR2X1 U77 ( .A(ab_27__1_), .B(ab_28__0_), .Y(SUMB_1__27_) );
  XOR2X1 U78 ( .A(ab_28__1_), .B(ab_29__0_), .Y(SUMB_1__28_) );
  XOR2X1 U79 ( .A(ab_29__1_), .B(ab_30__0_), .Y(SUMB_1__29_) );
  XOR2X1 U80 ( .A(CARRYB_30__0_), .B(SUMB_30__1_), .Y(PRODUCT[31]) );
  AND2X1 U81 ( .A(A[9]), .B(n48), .Y(ab_9__8_) );
  AND2X1 U82 ( .A(n46), .B(A[9]), .Y(ab_9__7_) );
  AND2X1 U83 ( .A(n46), .B(n48), .Y(ab_8__7_) );
  AND2X1 U84 ( .A(n44), .B(A[9]), .Y(ab_9__6_) );
  AND2X1 U85 ( .A(n44), .B(n48), .Y(ab_8__6_) );
  AND2X1 U86 ( .A(n44), .B(n46), .Y(ab_7__6_) );
  AND2X1 U87 ( .A(n42), .B(A[9]), .Y(ab_9__5_) );
  AND2X1 U88 ( .A(n42), .B(n48), .Y(ab_8__5_) );
  AND2X1 U89 ( .A(n42), .B(n46), .Y(ab_7__5_) );
  AND2X1 U90 ( .A(n42), .B(n44), .Y(ab_6__5_) );
  AND2X1 U91 ( .A(n40), .B(A[9]), .Y(ab_9__4_) );
  AND2X1 U92 ( .A(n40), .B(n48), .Y(ab_8__4_) );
  AND2X1 U93 ( .A(n40), .B(n46), .Y(ab_7__4_) );
  AND2X1 U94 ( .A(n40), .B(n44), .Y(ab_6__4_) );
  AND2X1 U95 ( .A(n40), .B(n42), .Y(ab_5__4_) );
  AND2X1 U96 ( .A(n38), .B(A[9]), .Y(ab_9__3_) );
  AND2X1 U97 ( .A(n38), .B(n48), .Y(ab_8__3_) );
  AND2X1 U98 ( .A(n38), .B(n46), .Y(ab_7__3_) );
  AND2X1 U99 ( .A(n38), .B(n44), .Y(ab_6__3_) );
  AND2X1 U100 ( .A(n38), .B(n42), .Y(ab_5__3_) );
  AND2X1 U101 ( .A(n38), .B(n40), .Y(ab_4__3_) );
  AND2X1 U102 ( .A(n36), .B(A[9]), .Y(ab_9__2_) );
  AND2X1 U103 ( .A(n36), .B(n48), .Y(ab_8__2_) );
  AND2X1 U104 ( .A(n36), .B(n46), .Y(ab_7__2_) );
  AND2X1 U105 ( .A(n36), .B(n44), .Y(ab_6__2_) );
  AND2X1 U106 ( .A(n36), .B(n42), .Y(ab_5__2_) );
  AND2X1 U107 ( .A(n36), .B(n40), .Y(ab_4__2_) );
  AND2X1 U108 ( .A(n36), .B(n38), .Y(ab_3__2_) );
  AND2X1 U109 ( .A(B[29]), .B(n36), .Y(ab_2__29_) );
  AND2X1 U110 ( .A(B[28]), .B(n38), .Y(ab_3__28_) );
  AND2X1 U111 ( .A(B[28]), .B(n36), .Y(ab_2__28_) );
  AND2X1 U112 ( .A(B[27]), .B(n40), .Y(ab_4__27_) );
  AND2X1 U113 ( .A(B[27]), .B(n38), .Y(ab_3__27_) );
  AND2X1 U114 ( .A(B[27]), .B(n36), .Y(ab_2__27_) );
  AND2X1 U115 ( .A(B[26]), .B(n42), .Y(ab_5__26_) );
  AND2X1 U116 ( .A(B[26]), .B(n40), .Y(ab_4__26_) );
  AND2X1 U117 ( .A(B[26]), .B(n38), .Y(ab_3__26_) );
  AND2X1 U118 ( .A(B[26]), .B(n36), .Y(ab_2__26_) );
  AND2X1 U119 ( .A(B[25]), .B(n44), .Y(ab_6__25_) );
  AND2X1 U120 ( .A(B[25]), .B(n42), .Y(ab_5__25_) );
  AND2X1 U121 ( .A(B[25]), .B(n40), .Y(ab_4__25_) );
  AND2X1 U122 ( .A(B[25]), .B(n38), .Y(ab_3__25_) );
  AND2X1 U123 ( .A(B[25]), .B(n36), .Y(ab_2__25_) );
  AND2X1 U124 ( .A(B[24]), .B(n46), .Y(ab_7__24_) );
  AND2X1 U125 ( .A(B[24]), .B(n44), .Y(ab_6__24_) );
  AND2X1 U126 ( .A(B[24]), .B(n42), .Y(ab_5__24_) );
  AND2X1 U127 ( .A(B[24]), .B(n40), .Y(ab_4__24_) );
  AND2X1 U128 ( .A(B[24]), .B(n38), .Y(ab_3__24_) );
  AND2X1 U129 ( .A(B[24]), .B(n36), .Y(ab_2__24_) );
  AND2X1 U130 ( .A(B[23]), .B(n48), .Y(ab_8__23_) );
  AND2X1 U131 ( .A(B[23]), .B(n46), .Y(ab_7__23_) );
  AND2X1 U132 ( .A(B[23]), .B(n44), .Y(ab_6__23_) );
  AND2X1 U133 ( .A(B[23]), .B(n42), .Y(ab_5__23_) );
  AND2X1 U134 ( .A(B[23]), .B(n40), .Y(ab_4__23_) );
  AND2X1 U135 ( .A(B[23]), .B(n38), .Y(ab_3__23_) );
  AND2X1 U136 ( .A(B[23]), .B(n36), .Y(ab_2__23_) );
  AND2X1 U137 ( .A(B[22]), .B(A[9]), .Y(ab_9__22_) );
  AND2X1 U138 ( .A(B[22]), .B(n48), .Y(ab_8__22_) );
  AND2X1 U139 ( .A(B[22]), .B(n46), .Y(ab_7__22_) );
  AND2X1 U140 ( .A(B[22]), .B(n44), .Y(ab_6__22_) );
  AND2X1 U141 ( .A(B[22]), .B(n42), .Y(ab_5__22_) );
  AND2X1 U142 ( .A(B[22]), .B(n40), .Y(ab_4__22_) );
  AND2X1 U143 ( .A(B[22]), .B(n38), .Y(ab_3__22_) );
  AND2X1 U144 ( .A(B[22]), .B(n36), .Y(ab_2__22_) );
  AND2X1 U145 ( .A(B[21]), .B(A[9]), .Y(ab_9__21_) );
  AND2X1 U146 ( .A(B[21]), .B(n48), .Y(ab_8__21_) );
  AND2X1 U147 ( .A(B[21]), .B(n46), .Y(ab_7__21_) );
  AND2X1 U148 ( .A(B[21]), .B(n44), .Y(ab_6__21_) );
  AND2X1 U149 ( .A(B[21]), .B(n42), .Y(ab_5__21_) );
  AND2X1 U150 ( .A(B[21]), .B(n40), .Y(ab_4__21_) );
  AND2X1 U151 ( .A(B[21]), .B(n38), .Y(ab_3__21_) );
  AND2X1 U152 ( .A(B[21]), .B(n36), .Y(ab_2__21_) );
  AND2X1 U153 ( .A(B[20]), .B(A[9]), .Y(ab_9__20_) );
  AND2X1 U154 ( .A(B[20]), .B(n48), .Y(ab_8__20_) );
  AND2X1 U155 ( .A(B[20]), .B(n46), .Y(ab_7__20_) );
  AND2X1 U156 ( .A(B[20]), .B(n44), .Y(ab_6__20_) );
  AND2X1 U157 ( .A(B[20]), .B(n42), .Y(ab_5__20_) );
  AND2X1 U158 ( .A(B[20]), .B(n40), .Y(ab_4__20_) );
  AND2X1 U159 ( .A(B[20]), .B(n38), .Y(ab_3__20_) );
  AND2X1 U160 ( .A(B[20]), .B(n36), .Y(ab_2__20_) );
  AND2X1 U161 ( .A(n34), .B(A[9]), .Y(ab_9__1_) );
  AND2X1 U162 ( .A(n34), .B(n48), .Y(ab_8__1_) );
  AND2X1 U163 ( .A(n34), .B(n46), .Y(ab_7__1_) );
  AND2X1 U164 ( .A(n34), .B(n44), .Y(ab_6__1_) );
  AND2X1 U165 ( .A(n34), .B(n42), .Y(ab_5__1_) );
  AND2X1 U166 ( .A(n34), .B(n40), .Y(ab_4__1_) );
  AND2X1 U167 ( .A(n34), .B(n38), .Y(ab_3__1_) );
  AND2X1 U168 ( .A(n34), .B(B[30]), .Y(ab_30__1_) );
  AND2X1 U169 ( .A(n34), .B(n36), .Y(ab_2__1_) );
  AND2X1 U170 ( .A(n34), .B(B[29]), .Y(ab_29__1_) );
  AND2X1 U171 ( .A(n34), .B(B[28]), .Y(ab_28__1_) );
  AND2X1 U172 ( .A(n34), .B(B[27]), .Y(ab_27__1_) );
  AND2X1 U173 ( .A(n34), .B(B[26]), .Y(ab_26__1_) );
  AND2X1 U174 ( .A(n34), .B(B[25]), .Y(ab_25__1_) );
  AND2X1 U175 ( .A(n34), .B(B[24]), .Y(ab_24__1_) );
  AND2X1 U176 ( .A(n34), .B(B[23]), .Y(ab_23__1_) );
  AND2X1 U177 ( .A(n34), .B(B[22]), .Y(ab_22__1_) );
  AND2X1 U178 ( .A(n34), .B(B[21]), .Y(ab_21__1_) );
  AND2X1 U179 ( .A(n34), .B(B[20]), .Y(ab_20__1_) );
  AND2X1 U180 ( .A(B[19]), .B(A[9]), .Y(ab_9__19_) );
  AND2X1 U181 ( .A(B[19]), .B(n48), .Y(ab_8__19_) );
  AND2X1 U182 ( .A(B[19]), .B(n46), .Y(ab_7__19_) );
  AND2X1 U183 ( .A(B[19]), .B(n44), .Y(ab_6__19_) );
  AND2X1 U184 ( .A(B[19]), .B(n42), .Y(ab_5__19_) );
  AND2X1 U185 ( .A(B[19]), .B(n40), .Y(ab_4__19_) );
  AND2X1 U186 ( .A(B[19]), .B(n38), .Y(ab_3__19_) );
  AND2X1 U187 ( .A(B[19]), .B(n36), .Y(ab_2__19_) );
  AND2X1 U188 ( .A(B[19]), .B(n34), .Y(ab_1__19_) );
  AND2X1 U189 ( .A(B[18]), .B(A[9]), .Y(ab_9__18_) );
  AND2X1 U190 ( .A(B[18]), .B(n48), .Y(ab_8__18_) );
  AND2X1 U191 ( .A(B[18]), .B(n46), .Y(ab_7__18_) );
  AND2X1 U192 ( .A(B[18]), .B(n44), .Y(ab_6__18_) );
  AND2X1 U193 ( .A(B[18]), .B(n42), .Y(ab_5__18_) );
  AND2X1 U194 ( .A(B[18]), .B(n40), .Y(ab_4__18_) );
  AND2X1 U195 ( .A(B[18]), .B(n38), .Y(ab_3__18_) );
  AND2X1 U196 ( .A(B[18]), .B(n36), .Y(ab_2__18_) );
  AND2X1 U197 ( .A(B[18]), .B(n34), .Y(ab_1__18_) );
  AND2X1 U198 ( .A(B[17]), .B(A[9]), .Y(ab_9__17_) );
  AND2X1 U199 ( .A(B[17]), .B(n48), .Y(ab_8__17_) );
  AND2X1 U200 ( .A(B[17]), .B(n46), .Y(ab_7__17_) );
  AND2X1 U201 ( .A(B[17]), .B(n44), .Y(ab_6__17_) );
  AND2X1 U202 ( .A(B[17]), .B(n42), .Y(ab_5__17_) );
  AND2X1 U203 ( .A(B[17]), .B(n40), .Y(ab_4__17_) );
  AND2X1 U204 ( .A(B[17]), .B(n38), .Y(ab_3__17_) );
  AND2X1 U205 ( .A(B[17]), .B(n36), .Y(ab_2__17_) );
  AND2X1 U206 ( .A(B[17]), .B(n34), .Y(ab_1__17_) );
  AND2X1 U207 ( .A(B[16]), .B(A[9]), .Y(ab_9__16_) );
  AND2X1 U208 ( .A(B[16]), .B(n48), .Y(ab_8__16_) );
  AND2X1 U209 ( .A(B[16]), .B(n46), .Y(ab_7__16_) );
  AND2X1 U210 ( .A(B[16]), .B(n44), .Y(ab_6__16_) );
  AND2X1 U211 ( .A(B[16]), .B(n42), .Y(ab_5__16_) );
  AND2X1 U212 ( .A(B[16]), .B(n40), .Y(ab_4__16_) );
  AND2X1 U213 ( .A(B[16]), .B(n38), .Y(ab_3__16_) );
  AND2X1 U214 ( .A(B[16]), .B(n36), .Y(ab_2__16_) );
  AND2X1 U215 ( .A(B[16]), .B(n34), .Y(ab_1__16_) );
  AND2X1 U216 ( .A(B[15]), .B(A[9]), .Y(ab_9__15_) );
  AND2X1 U217 ( .A(B[15]), .B(n48), .Y(ab_8__15_) );
  AND2X1 U218 ( .A(B[15]), .B(n46), .Y(ab_7__15_) );
  AND2X1 U219 ( .A(B[15]), .B(n44), .Y(ab_6__15_) );
  AND2X1 U220 ( .A(B[15]), .B(n42), .Y(ab_5__15_) );
  AND2X1 U221 ( .A(B[15]), .B(n40), .Y(ab_4__15_) );
  AND2X1 U222 ( .A(B[15]), .B(n38), .Y(ab_3__15_) );
  AND2X1 U223 ( .A(B[15]), .B(n36), .Y(ab_2__15_) );
  AND2X1 U224 ( .A(B[15]), .B(n34), .Y(ab_1__15_) );
  AND2X1 U225 ( .A(B[15]), .B(B[16]), .Y(ab_16__15_) );
  AND2X1 U226 ( .A(B[14]), .B(A[9]), .Y(ab_9__14_) );
  AND2X1 U227 ( .A(B[14]), .B(n48), .Y(ab_8__14_) );
  AND2X1 U228 ( .A(B[14]), .B(n46), .Y(ab_7__14_) );
  AND2X1 U229 ( .A(B[14]), .B(n44), .Y(ab_6__14_) );
  AND2X1 U230 ( .A(B[14]), .B(n42), .Y(ab_5__14_) );
  AND2X1 U231 ( .A(B[14]), .B(n40), .Y(ab_4__14_) );
  AND2X1 U232 ( .A(B[14]), .B(n38), .Y(ab_3__14_) );
  AND2X1 U233 ( .A(B[14]), .B(n36), .Y(ab_2__14_) );
  AND2X1 U234 ( .A(B[14]), .B(n34), .Y(ab_1__14_) );
  AND2X1 U235 ( .A(B[14]), .B(B[17]), .Y(ab_17__14_) );
  AND2X1 U236 ( .A(B[14]), .B(B[16]), .Y(ab_16__14_) );
  AND2X1 U237 ( .A(B[14]), .B(B[15]), .Y(ab_15__14_) );
  AND2X1 U238 ( .A(B[13]), .B(A[9]), .Y(ab_9__13_) );
  AND2X1 U239 ( .A(B[13]), .B(n48), .Y(ab_8__13_) );
  AND2X1 U240 ( .A(B[13]), .B(n46), .Y(ab_7__13_) );
  AND2X1 U241 ( .A(B[13]), .B(n44), .Y(ab_6__13_) );
  AND2X1 U242 ( .A(B[13]), .B(n42), .Y(ab_5__13_) );
  AND2X1 U243 ( .A(B[13]), .B(n40), .Y(ab_4__13_) );
  AND2X1 U244 ( .A(B[13]), .B(n38), .Y(ab_3__13_) );
  AND2X1 U245 ( .A(B[13]), .B(n36), .Y(ab_2__13_) );
  AND2X1 U246 ( .A(B[13]), .B(n34), .Y(ab_1__13_) );
  AND2X1 U247 ( .A(B[13]), .B(B[18]), .Y(ab_18__13_) );
  AND2X1 U248 ( .A(B[13]), .B(B[17]), .Y(ab_17__13_) );
  AND2X1 U249 ( .A(B[13]), .B(B[16]), .Y(ab_16__13_) );
  AND2X1 U250 ( .A(B[13]), .B(B[15]), .Y(ab_15__13_) );
  AND2X1 U251 ( .A(B[13]), .B(B[14]), .Y(ab_14__13_) );
  AND2X1 U252 ( .A(A[12]), .B(A[9]), .Y(ab_9__12_) );
  AND2X1 U253 ( .A(A[12]), .B(n48), .Y(ab_8__12_) );
  AND2X1 U254 ( .A(A[12]), .B(n46), .Y(ab_7__12_) );
  AND2X1 U255 ( .A(A[12]), .B(n44), .Y(ab_6__12_) );
  AND2X1 U256 ( .A(A[12]), .B(n42), .Y(ab_5__12_) );
  AND2X1 U257 ( .A(A[12]), .B(n40), .Y(ab_4__12_) );
  AND2X1 U258 ( .A(A[12]), .B(n38), .Y(ab_3__12_) );
  AND2X1 U259 ( .A(A[12]), .B(n36), .Y(ab_2__12_) );
  AND2X1 U260 ( .A(A[12]), .B(n34), .Y(ab_1__12_) );
  AND2X1 U261 ( .A(A[12]), .B(B[19]), .Y(ab_19__12_) );
  AND2X1 U262 ( .A(A[12]), .B(B[18]), .Y(ab_18__12_) );
  AND2X1 U263 ( .A(A[12]), .B(B[17]), .Y(ab_17__12_) );
  AND2X1 U264 ( .A(A[12]), .B(B[16]), .Y(ab_16__12_) );
  AND2X1 U265 ( .A(A[12]), .B(B[15]), .Y(ab_15__12_) );
  AND2X1 U266 ( .A(A[12]), .B(B[14]), .Y(ab_14__12_) );
  AND2X1 U267 ( .A(A[12]), .B(B[13]), .Y(ab_13__12_) );
  AND2X1 U268 ( .A(n52), .B(A[9]), .Y(ab_9__11_) );
  AND2X1 U269 ( .A(n52), .B(n48), .Y(ab_8__11_) );
  AND2X1 U270 ( .A(n52), .B(n46), .Y(ab_7__11_) );
  AND2X1 U271 ( .A(n52), .B(n44), .Y(ab_6__11_) );
  AND2X1 U272 ( .A(n52), .B(n42), .Y(ab_5__11_) );
  AND2X1 U273 ( .A(n52), .B(n40), .Y(ab_4__11_) );
  AND2X1 U274 ( .A(n52), .B(n38), .Y(ab_3__11_) );
  AND2X1 U275 ( .A(n52), .B(n36), .Y(ab_2__11_) );
  AND2X1 U276 ( .A(n52), .B(B[20]), .Y(ab_20__11_) );
  AND2X1 U277 ( .A(n52), .B(n34), .Y(ab_1__11_) );
  AND2X1 U278 ( .A(n52), .B(B[19]), .Y(ab_19__11_) );
  AND2X1 U279 ( .A(n52), .B(B[18]), .Y(ab_18__11_) );
  AND2X1 U280 ( .A(n52), .B(B[17]), .Y(ab_17__11_) );
  AND2X1 U281 ( .A(n52), .B(B[16]), .Y(ab_16__11_) );
  AND2X1 U282 ( .A(n52), .B(B[15]), .Y(ab_15__11_) );
  AND2X1 U283 ( .A(n52), .B(B[14]), .Y(ab_14__11_) );
  AND2X1 U284 ( .A(n52), .B(B[13]), .Y(ab_13__11_) );
  AND2X1 U285 ( .A(n52), .B(A[12]), .Y(ab_12__11_) );
  AND2X1 U286 ( .A(n50), .B(A[9]), .Y(ab_9__10_) );
  AND2X1 U287 ( .A(n50), .B(n48), .Y(ab_8__10_) );
  AND2X1 U288 ( .A(n50), .B(n46), .Y(ab_7__10_) );
  AND2X1 U289 ( .A(n50), .B(n44), .Y(ab_6__10_) );
  AND2X1 U290 ( .A(n50), .B(n42), .Y(ab_5__10_) );
  AND2X1 U291 ( .A(n50), .B(n40), .Y(ab_4__10_) );
  AND2X1 U292 ( .A(n50), .B(n38), .Y(ab_3__10_) );
  AND2X1 U293 ( .A(n50), .B(n36), .Y(ab_2__10_) );
  AND2X1 U294 ( .A(n50), .B(B[21]), .Y(ab_21__10_) );
  AND2X1 U295 ( .A(n50), .B(B[20]), .Y(ab_20__10_) );
  AND2X1 U296 ( .A(n50), .B(n34), .Y(ab_1__10_) );
  AND2X1 U297 ( .A(n50), .B(B[19]), .Y(ab_19__10_) );
  AND2X1 U298 ( .A(n50), .B(B[18]), .Y(ab_18__10_) );
  AND2X1 U299 ( .A(n50), .B(B[17]), .Y(ab_17__10_) );
  AND2X1 U300 ( .A(n50), .B(B[16]), .Y(ab_16__10_) );
  AND2X1 U301 ( .A(n50), .B(B[15]), .Y(ab_15__10_) );
  AND2X1 U302 ( .A(n50), .B(B[14]), .Y(ab_14__10_) );
  AND2X1 U303 ( .A(n50), .B(B[13]), .Y(ab_13__10_) );
  AND2X1 U304 ( .A(n50), .B(A[12]), .Y(ab_12__10_) );
  AND2X1 U305 ( .A(n50), .B(n52), .Y(ab_11__10_) );
  AND2X1 U306 ( .A(B[0]), .B(B[9]), .Y(ab_9__0_) );
  AND2X1 U307 ( .A(B[0]), .B(n48), .Y(ab_8__0_) );
  AND2X1 U308 ( .A(B[0]), .B(n46), .Y(ab_7__0_) );
  AND2X1 U309 ( .A(B[0]), .B(n44), .Y(ab_6__0_) );
  AND2X1 U310 ( .A(B[0]), .B(n42), .Y(ab_5__0_) );
  AND2X1 U311 ( .A(B[0]), .B(n40), .Y(ab_4__0_) );
  AND2X1 U312 ( .A(B[0]), .B(n38), .Y(ab_3__0_) );
  AND2X1 U313 ( .A(B[0]), .B(B[30]), .Y(ab_30__0_) );
  AND2X1 U314 ( .A(B[0]), .B(n36), .Y(ab_2__0_) );
  AND2X1 U315 ( .A(B[0]), .B(B[29]), .Y(ab_29__0_) );
  AND2X1 U316 ( .A(B[0]), .B(B[28]), .Y(ab_28__0_) );
  AND2X1 U317 ( .A(B[0]), .B(B[27]), .Y(ab_27__0_) );
  AND2X1 U318 ( .A(B[0]), .B(B[26]), .Y(ab_26__0_) );
  AND2X1 U319 ( .A(B[0]), .B(B[25]), .Y(ab_25__0_) );
  AND2X1 U320 ( .A(B[0]), .B(B[24]), .Y(ab_24__0_) );
  AND2X1 U321 ( .A(B[0]), .B(B[23]), .Y(ab_23__0_) );
  AND2X1 U322 ( .A(B[0]), .B(B[22]), .Y(ab_22__0_) );
  AND2X1 U323 ( .A(B[0]), .B(B[21]), .Y(ab_21__0_) );
  AND2X1 U324 ( .A(B[0]), .B(B[20]), .Y(ab_20__0_) );
  AND2X1 U325 ( .A(B[0]), .B(B[19]), .Y(ab_19__0_) );
  AND2X1 U326 ( .A(B[0]), .B(B[18]), .Y(ab_18__0_) );
  AND2X1 U327 ( .A(B[0]), .B(B[17]), .Y(ab_17__0_) );
  AND2X1 U328 ( .A(B[0]), .B(B[16]), .Y(ab_16__0_) );
  AND2X1 U329 ( .A(B[0]), .B(B[15]), .Y(ab_15__0_) );
  AND2X1 U330 ( .A(B[0]), .B(B[14]), .Y(ab_14__0_) );
  AND2X1 U331 ( .A(B[0]), .B(B[13]), .Y(ab_13__0_) );
  AND2X1 U332 ( .A(B[0]), .B(B[12]), .Y(ab_12__0_) );
  AND2X1 U333 ( .A(B[0]), .B(n52), .Y(ab_11__0_) );
  AND2X1 U334 ( .A(B[0]), .B(n50), .Y(ab_10__0_) );
  AND2X1 U335 ( .A(n34), .B(B[0]), .Y(CARRYB_1__0_) );
endmodule


module square_root_finder_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_, ab_28__3_,
         ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_, ab_27__2_,
         ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_, ab_26__2_,
         ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_, ab_25__3_,
         ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_, ab_24__5_,
         ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_, ab_22__6_,
         ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_, ab_22__0_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__11_,
         ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_, ab_20__5_,
         ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_, ab_19__12_,
         ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_, ab_19__6_,
         ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_, ab_19__0_,
         ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_, ab_18__8_,
         ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_, ab_18__2_,
         ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__15_,
         ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_,
         ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_,
         ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_, ab_15__14_, ab_15__13_,
         ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_,
         ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_,
         ab_15__0_, ab_14__17_, ab_14__16_, ab_14__15_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_,
         ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_,
         ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_, ab_12__15_,
         ab_12__14_, ab_12__13_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_,
         ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_,
         ab_12__1_, ab_12__0_, ab_11__20_, ab_11__19_, ab_11__18_, ab_11__17_,
         ab_11__16_, ab_11__15_, ab_11__14_, ab_11__13_, ab_11__12_,
         ab_11__10_, ab_11__9_, ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_,
         ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_,
         ab_10__20_, ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_,
         ab_10__15_, ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_,
         ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_,
         ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__6_, ab_7__5_,
         ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__26_,
         ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_, ab_5__20_,
         ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_, ab_5__14_,
         ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_, ab_5__8_,
         ab_5__7_, ab_5__6_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_,
         ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__28_, ab_3__27_, ab_3__26_, ab_3__25_,
         ab_3__24_, ab_3__23_, ab_3__22_, ab_3__21_, ab_3__20_, ab_3__19_,
         ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_, ab_3__14_, ab_3__13_,
         ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_, ab_3__8_, ab_3__7_,
         ab_3__6_, ab_3__5_, ab_3__4_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_,
         ab_2__28_, ab_2__27_, ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_,
         ab_2__22_, ab_2__21_, ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_,
         ab_2__16_, ab_2__15_, ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_,
         ab_2__10_, ab_2__9_, ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_,
         ab_1__27_, ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_,
         ab_1__21_, ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_,
         ab_1__15_, ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_,
         ab_1__9_, ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_,
         ab_1__2_, ab_1__0_, ab_0__30_, ab_0__29_, ab_0__28_, ab_0__27_,
         ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_, ab_0__21_,
         ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_, ab_0__15_,
         ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_, ab_0__9_,
         ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_,
         ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_15__16_, SUMB_15__15_,
         SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_, SUMB_15__10_,
         SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__17_,
         SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_, SUMB_14__12_,
         SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_, SUMB_14__7_,
         SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_,
         SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_,
         SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_,
         SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_,
         SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__19_,
         SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_, SUMB_12__14_,
         SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_, SUMB_12__9_,
         SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_,
         SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_, SUMB_10__20_,
         SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_, SUMB_10__15_,
         SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_, SUMB_10__10_,
         SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__22_,
         SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_, SUMB_9__17_,
         SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_, SUMB_9__12_,
         SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_, SUMB_9__7_,
         SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_,
         SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_,
         SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_,
         SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_,
         SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_,
         SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__24_,
         SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_, SUMB_7__19_,
         SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_, SUMB_7__14_,
         SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_, SUMB_7__9_,
         SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_,
         SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_, SUMB_6__24_,
         SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_, SUMB_5__25_,
         SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_, SUMB_5__20_,
         SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_, SUMB_5__15_,
         SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_, SUMB_5__10_,
         SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__27_,
         SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_, SUMB_4__22_,
         SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_, SUMB_4__17_,
         SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_, SUMB_4__12_,
         SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_, SUMB_4__7_,
         SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_,
         SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_, SUMB_3__25_,
         SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_,
         SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_,
         SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_,
         SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_,
         SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__29_,
         SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_, SUMB_2__24_,
         SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_, SUMB_2__19_,
         SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_, SUMB_2__14_,
         SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_, SUMB_2__9_,
         SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_,
         SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__29_, SUMB_1__28_,
         SUMB_1__27_, SUMB_1__26_, SUMB_1__25_, SUMB_1__24_, SUMB_1__23_,
         SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_, SUMB_1__18_,
         SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_, SUMB_1__13_,
         SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_, SUMB_1__8_,
         SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_, CARRYB_29__1_, CARRYB_29__0_,
         CARRYB_28__2_, CARRYB_28__1_, CARRYB_28__0_, CARRYB_27__3_,
         CARRYB_27__2_, CARRYB_27__1_, CARRYB_27__0_, CARRYB_26__4_,
         CARRYB_26__3_, CARRYB_26__2_, CARRYB_26__1_, CARRYB_26__0_,
         CARRYB_25__5_, CARRYB_25__4_, CARRYB_25__3_, CARRYB_25__2_,
         CARRYB_25__1_, CARRYB_25__0_, CARRYB_24__6_, CARRYB_24__5_,
         CARRYB_24__4_, CARRYB_24__3_, CARRYB_24__2_, CARRYB_24__1_,
         CARRYB_24__0_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__8_, CARRYB_22__7_, CARRYB_22__6_,
         CARRYB_22__5_, CARRYB_22__4_, CARRYB_22__3_, CARRYB_22__2_,
         CARRYB_22__1_, CARRYB_22__0_, CARRYB_21__9_, CARRYB_21__8_,
         CARRYB_21__7_, CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_,
         CARRYB_21__3_, CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_,
         CARRYB_20__10_, CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_,
         CARRYB_20__6_, CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_,
         CARRYB_20__2_, CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__11_,
         CARRYB_19__10_, CARRYB_19__9_, CARRYB_19__8_, CARRYB_19__7_,
         CARRYB_19__6_, CARRYB_19__5_, CARRYB_19__4_, CARRYB_19__3_,
         CARRYB_19__2_, CARRYB_19__1_, CARRYB_19__0_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_, CARRYB_17__10_,
         CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_, CARRYB_17__6_,
         CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_, CARRYB_17__2_,
         CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__14_, CARRYB_16__13_,
         CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_, CARRYB_16__9_,
         CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_, CARRYB_16__5_,
         CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_,
         CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_, SUMB_29__1_, SUMB_28__3_,
         SUMB_28__2_, SUMB_28__1_, SUMB_27__4_, SUMB_27__3_, SUMB_27__2_,
         SUMB_27__1_, SUMB_26__5_, SUMB_26__4_, SUMB_26__3_, SUMB_26__2_,
         SUMB_26__1_, SUMB_25__6_, SUMB_25__5_, SUMB_25__4_, SUMB_25__3_,
         SUMB_25__2_, SUMB_25__1_, SUMB_24__7_, SUMB_24__6_, SUMB_24__5_,
         SUMB_24__4_, SUMB_24__3_, SUMB_24__2_, SUMB_24__1_, SUMB_23__8_,
         SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_, SUMB_23__3_,
         SUMB_23__2_, SUMB_23__1_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__10_, SUMB_21__9_, SUMB_21__8_, SUMB_21__7_,
         SUMB_21__6_, SUMB_21__5_, SUMB_21__4_, SUMB_21__3_, SUMB_21__2_,
         SUMB_21__1_, SUMB_20__11_, SUMB_20__10_, SUMB_20__9_, SUMB_20__8_,
         SUMB_20__7_, SUMB_20__6_, SUMB_20__5_, SUMB_20__4_, SUMB_20__3_,
         SUMB_20__2_, SUMB_20__1_, SUMB_19__12_, SUMB_19__11_, SUMB_19__10_,
         SUMB_19__9_, SUMB_19__8_, SUMB_19__7_, SUMB_19__6_, SUMB_19__5_,
         SUMB_19__4_, SUMB_19__3_, SUMB_19__2_, SUMB_19__1_, SUMB_18__13_,
         SUMB_18__12_, SUMB_18__11_, SUMB_18__10_, SUMB_18__9_, SUMB_18__8_,
         SUMB_18__7_, SUMB_18__6_, SUMB_18__5_, SUMB_18__4_, SUMB_18__3_,
         SUMB_18__2_, SUMB_18__1_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__15_, SUMB_16__14_, SUMB_16__13_, SUMB_16__12_,
         SUMB_16__11_, SUMB_16__10_, SUMB_16__9_, SUMB_16__8_, SUMB_16__7_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89;

  ADDFX2 S2_2_28 ( .A(ab_2__28_), .B(n35), .CI(SUMB_1__29_), .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  ADDFX2 S2_2_27 ( .A(ab_2__27_), .B(n34), .CI(SUMB_1__28_), .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  ADDFX2 S2_2_26 ( .A(ab_2__26_), .B(n33), .CI(SUMB_1__27_), .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  ADDFX2 S2_2_25 ( .A(ab_2__25_), .B(n32), .CI(SUMB_1__26_), .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  ADDFX2 S2_2_24 ( .A(ab_2__24_), .B(n31), .CI(SUMB_1__25_), .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  ADDFX2 S2_2_23 ( .A(ab_2__23_), .B(n30), .CI(SUMB_1__24_), .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  ADDFX2 S2_2_22 ( .A(ab_2__22_), .B(n29), .CI(SUMB_1__23_), .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  ADDFX2 S2_2_21 ( .A(ab_2__21_), .B(n28), .CI(SUMB_1__22_), .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  ADDFX2 S2_2_20 ( .A(ab_2__20_), .B(n27), .CI(SUMB_1__21_), .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  ADDFX2 S2_2_19 ( .A(ab_2__19_), .B(n26), .CI(SUMB_1__20_), .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  ADDFX2 S2_2_18 ( .A(ab_2__18_), .B(n25), .CI(SUMB_1__19_), .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  ADDFX2 S2_2_17 ( .A(ab_2__17_), .B(n24), .CI(SUMB_1__18_), .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  ADDFX2 S2_2_16 ( .A(ab_2__16_), .B(n23), .CI(SUMB_1__17_), .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  XOR3X2 S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .C(SUMB_22__9_), .Y(
        SUMB_23__8_) );
  XOR3X2 S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .C(SUMB_23__8_), .Y(
        SUMB_24__7_) );
  XOR3X2 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .C(SUMB_20__11_), .Y(
        SUMB_21__10_) );
  XOR3X2 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .C(SUMB_21__10_), .Y(
        SUMB_22__9_) );
  XOR3X2 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .C(SUMB_18__13_), .Y(
        SUMB_19__12_) );
  XOR3X2 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .C(SUMB_19__12_), .Y(
        SUMB_20__11_) );
  XOR3X2 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .C(SUMB_16__15_), .Y(
        SUMB_17__14_) );
  XOR3X2 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .C(SUMB_17__14_), .Y(
        SUMB_18__13_) );
  XOR3X2 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .C(SUMB_14__17_), .Y(
        SUMB_15__16_) );
  XOR3X2 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .C(SUMB_15__16_), .Y(
        SUMB_16__15_) );
  XOR3X2 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .C(SUMB_12__19_), .Y(
        SUMB_13__18_) );
  XOR3X2 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .C(SUMB_13__18_), .Y(
        SUMB_14__17_) );
  XOR3X2 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .C(SUMB_10__21_), .Y(
        SUMB_11__20_) );
  XOR3X2 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .C(SUMB_11__20_), .Y(
        SUMB_12__19_) );
  XOR3X2 S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .C(SUMB_8__23_), .Y(
        SUMB_9__22_) );
  XOR3X2 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .C(SUMB_9__22_), .Y(
        SUMB_10__21_) );
  XOR3X2 S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .C(SUMB_6__25_), .Y(
        SUMB_7__24_) );
  XOR3X2 S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .C(SUMB_7__24_), .Y(
        SUMB_8__23_) );
  XOR3X2 S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .C(SUMB_4__27_), .Y(
        SUMB_5__26_) );
  XOR3X2 S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .C(SUMB_5__26_), .Y(
        SUMB_6__25_) );
  XOR3X2 S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .C(SUMB_2__29_), .Y(
        SUMB_3__28_) );
  XOR3X2 S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .C(SUMB_3__28_), .Y(
        SUMB_4__27_) );
  XOR3X2 S2_2_29 ( .A(ab_2__29_), .B(n36), .C(ab_1__30_), .Y(SUMB_2__29_) );
  ADDFX2 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  ADDFX2 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  ADDFX2 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  ADDFX2 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  ADDFX2 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  ADDFX2 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  ADDFX2 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  ADDFX2 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  ADDFX2 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  ADDFX2 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  ADDFX2 S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  ADDFX2 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  ADDFX2 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  ADDFX2 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  ADDFX2 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  ADDFX2 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  ADDFX2 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  ADDFX2 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  ADDFX2 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  ADDFX2 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  ADDFX2 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  ADDFX2 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  ADDFX2 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  ADDFX2 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  ADDFX2 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  ADDFX2 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  ADDFX2 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  ADDFX2 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  ADDFX2 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  ADDFX2 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  ADDFX2 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  ADDFX2 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  ADDFX2 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  ADDFX2 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  ADDFX2 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  ADDFX2 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  ADDFX2 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  ADDFX2 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  ADDFX2 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  ADDFX2 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  ADDFX2 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  ADDFX2 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  ADDFX2 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  ADDFX2 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  ADDFX2 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  ADDFX2 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  ADDFX2 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  ADDFX2 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  ADDFX2 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  ADDFX2 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  ADDFX2 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  ADDFX2 S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  ADDFX2 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  ADDFX2 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  ADDFX2 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  ADDFX2 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  ADDFX2 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  ADDFX2 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  ADDFX2 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  ADDFX2 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  ADDFX2 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  ADDFX2 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  ADDFX2 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFX2 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  ADDFX2 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  ADDFX2 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  ADDFX2 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  ADDFX2 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  ADDFX2 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  ADDFX2 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  ADDFX2 S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), .CO(
        CARRYB_7__23_), .S(SUMB_7__23_) );
  ADDFX2 S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  ADDFX2 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  ADDFX2 S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), .CO(
        CARRYB_6__23_), .S(SUMB_6__23_) );
  ADDFX2 S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  ADDFX2 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  ADDFX2 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  ADDFX2 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  ADDFX2 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  ADDFX2 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  ADDFX2 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  ADDFX2 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  ADDFX2 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  ADDFX2 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  ADDFX2 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  ADDFX2 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  ADDFX2 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  ADDFX2 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  ADDFX2 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  ADDFX2 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  ADDFX2 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  ADDFX2 S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), .CO(
        CARRYB_24__6_), .S(SUMB_24__6_) );
  ADDFX2 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  ADDFX2 S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), .CO(
        CARRYB_4__26_), .S(SUMB_4__26_) );
  ADDFX2 S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), .CO(
        CARRYB_4__25_), .S(SUMB_4__25_) );
  ADDFX2 S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), .CO(
        CARRYB_4__24_), .S(SUMB_4__24_) );
  ADDFX2 S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), .CO(
        CARRYB_4__23_), .S(SUMB_4__23_) );
  ADDFX2 S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  ADDFX2 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  ADDFX2 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  ADDFX2 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  ADDFX2 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  ADDFX2 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  ADDFX2 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  ADDFX2 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  ADDFX2 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  ADDFX2 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  ADDFX2 S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  ADDFX2 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  ADDFX2 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  ADDFX2 S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), .CO(
        CARRYB_6__24_), .S(SUMB_6__24_) );
  ADDFX2 S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), .CO(
        CARRYB_5__25_), .S(SUMB_5__25_) );
  ADDFX2 S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), .CO(
        CARRYB_5__24_), .S(SUMB_5__24_) );
  ADDFX2 S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), .CO(
        CARRYB_5__23_), .S(SUMB_5__23_) );
  ADDFX2 S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  ADDFX2 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  ADDFX2 S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), .CO(
        CARRYB_3__27_), .S(SUMB_3__27_) );
  ADDFX2 S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), .CO(
        CARRYB_3__26_), .S(SUMB_3__26_) );
  ADDFX2 S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), .CO(
        CARRYB_3__25_), .S(SUMB_3__25_) );
  ADDFX2 S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), .CO(
        CARRYB_3__24_), .S(SUMB_3__24_) );
  ADDFX2 S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), .CO(
        CARRYB_3__23_), .S(SUMB_3__23_) );
  ADDFX2 S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  ADDFX2 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  ADDFX2 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  ADDFX2 S2_12_12 ( .A(B[12]), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  ADDFX2 S2_15_15 ( .A(B[15]), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  ADDFX2 S2_14_14 ( .A(B[14]), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  ADDFX2 S2_13_13 ( .A(B[13]), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  ADDFX2 S2_11_11 ( .A(B[11]), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  ADDFX2 S2_10_10 ( .A(B[10]), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  ADDFX2 S2_9_9 ( .A(B[9]), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  ADDFX2 S2_8_8 ( .A(B[8]), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  ADDFX2 S2_7_7 ( .A(B[7]), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  ADDFX2 S2_6_6 ( .A(B[6]), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  XOR3X2 S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .C(SUMB_26__5_), .Y(
        SUMB_27__4_) );
  XOR3X2 S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .C(SUMB_27__4_), .Y(
        SUMB_28__3_) );
  XOR3X2 S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .C(SUMB_24__7_), .Y(
        SUMB_25__6_) );
  XOR3X2 S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .C(SUMB_25__6_), .Y(
        SUMB_26__5_) );
  ADDFX2 S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), .CO(
        CARRYB_30__0_), .S(PRODUCT[30]) );
  XOR3X2 S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .C(SUMB_28__3_), .Y(
        SUMB_29__2_) );
  XOR3X2 S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .C(SUMB_29__2_), .Y(
        SUMB_30__1_) );
  ADDFX2 S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), .CO(
        CARRYB_29__1_), .S(SUMB_29__1_) );
  ADDFX2 S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), .CO(
        CARRYB_29__0_), .S(PRODUCT[29]) );
  ADDFX2 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  ADDFX2 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  ADDFX2 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  ADDFX2 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  ADDFX2 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  ADDFX2 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(PRODUCT[19]) );
  ADDFX2 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  ADDFX2 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  ADDFX2 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  ADDFX2 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  ADDFX2 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  ADDFX2 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(PRODUCT[18]) );
  ADDFX2 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  ADDFX2 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  ADDFX2 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  ADDFX2 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  ADDFX2 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  ADDFX2 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(PRODUCT[17]) );
  ADDFX2 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFX2 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFX2 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFX2 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFX2 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFX2 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(PRODUCT[16]) );
  ADDFX2 S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), .CO(
        CARRYB_28__2_), .S(SUMB_28__2_) );
  ADDFX2 S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), .CO(
        CARRYB_28__1_), .S(SUMB_28__1_) );
  ADDFX2 S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), .CO(
        CARRYB_28__0_), .S(PRODUCT[28]) );
  ADDFX2 S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), .CO(
        CARRYB_27__3_), .S(SUMB_27__3_) );
  ADDFX2 S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), .CO(
        CARRYB_27__2_), .S(SUMB_27__2_) );
  ADDFX2 S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), .CO(
        CARRYB_27__1_), .S(SUMB_27__1_) );
  ADDFX2 S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), .CO(
        CARRYB_27__0_), .S(PRODUCT[27]) );
  ADDFX2 S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), .CO(
        CARRYB_26__4_), .S(SUMB_26__4_) );
  ADDFX2 S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), .CO(
        CARRYB_26__3_), .S(SUMB_26__3_) );
  ADDFX2 S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), .CO(
        CARRYB_26__2_), .S(SUMB_26__2_) );
  ADDFX2 S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), .CO(
        CARRYB_26__1_), .S(SUMB_26__1_) );
  ADDFX2 S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), .CO(
        CARRYB_26__0_), .S(PRODUCT[26]) );
  ADDFX2 S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), .CO(
        CARRYB_25__5_), .S(SUMB_25__5_) );
  ADDFX2 S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), .CO(
        CARRYB_25__4_), .S(SUMB_25__4_) );
  ADDFX2 S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), .CO(
        CARRYB_25__3_), .S(SUMB_25__3_) );
  ADDFX2 S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), .CO(
        CARRYB_25__2_), .S(SUMB_25__2_) );
  ADDFX2 S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), .CO(
        CARRYB_25__1_), .S(SUMB_25__1_) );
  ADDFX2 S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), .CO(
        CARRYB_25__0_), .S(PRODUCT[25]) );
  ADDFX2 S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), .CO(
        CARRYB_24__5_), .S(SUMB_24__5_) );
  ADDFX2 S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), .CO(
        CARRYB_24__4_), .S(SUMB_24__4_) );
  ADDFX2 S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), .CO(
        CARRYB_24__3_), .S(SUMB_24__3_) );
  ADDFX2 S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), .CO(
        CARRYB_24__2_), .S(SUMB_24__2_) );
  ADDFX2 S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), .CO(
        CARRYB_24__1_), .S(SUMB_24__1_) );
  ADDFX2 S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), .CO(
        CARRYB_24__0_), .S(PRODUCT[24]) );
  ADDFX2 S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  ADDFX2 S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  ADDFX2 S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  ADDFX2 S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  ADDFX2 S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  ADDFX2 S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(PRODUCT[23]) );
  ADDFX2 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  ADDFX2 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  ADDFX2 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  ADDFX2 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  ADDFX2 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  ADDFX2 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(PRODUCT[22]) );
  ADDFX2 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  ADDFX2 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  ADDFX2 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  ADDFX2 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  ADDFX2 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  ADDFX2 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(PRODUCT[21]) );
  ADDFX2 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  ADDFX2 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  ADDFX2 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  ADDFX2 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  ADDFX2 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  ADDFX2 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(PRODUCT[20]) );
  ADDFX2 S2_5_5 ( .A(B[5]), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  ADDFX2 S2_2_14 ( .A(ab_2__14_), .B(n22), .CI(SUMB_1__15_), .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  ADDFX2 S2_2_13 ( .A(ab_2__13_), .B(n21), .CI(SUMB_1__14_), .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  ADDFX2 S2_2_12 ( .A(ab_2__12_), .B(n20), .CI(SUMB_1__13_), .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  ADDFX2 S2_2_11 ( .A(ab_2__11_), .B(n17), .CI(SUMB_1__12_), .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  ADDFX2 S2_2_10 ( .A(ab_2__10_), .B(n16), .CI(SUMB_1__11_), .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  ADDFX2 S2_2_9 ( .A(ab_2__9_), .B(n15), .CI(SUMB_1__10_), .CO(CARRYB_2__9_), 
        .S(SUMB_2__9_) );
  ADDFX2 S2_2_8 ( .A(ab_2__8_), .B(n18), .CI(SUMB_1__9_), .CO(CARRYB_2__8_), 
        .S(SUMB_2__8_) );
  ADDFX2 S2_2_7 ( .A(ab_2__7_), .B(n14), .CI(SUMB_1__8_), .CO(CARRYB_2__7_), 
        .S(SUMB_2__7_) );
  ADDFX2 S2_2_6 ( .A(ab_2__6_), .B(n11), .CI(SUMB_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFX2 S2_2_15 ( .A(ab_2__15_), .B(n19), .CI(SUMB_1__16_), .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  ADDFX2 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  ADDFX2 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  ADDFX2 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  ADDFX2 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  ADDFX2 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  ADDFX2 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  ADDFX2 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  ADDFX2 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  ADDFX2 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  ADDFX2 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  ADDFX2 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  ADDFX2 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFX2 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  ADDFX2 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  ADDFX2 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  ADDFX2 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  ADDFX2 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  ADDFX2 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  ADDFX2 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  ADDFX2 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFX2 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  ADDFX2 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  ADDFX2 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  ADDFX2 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  ADDFX2 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  ADDFX2 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  ADDFX2 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  ADDFX2 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  ADDFX2 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFX2 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  ADDFX2 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  ADDFX2 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  ADDFX2 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  ADDFX2 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  ADDFX2 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  ADDFX2 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  ADDFX2 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  ADDFX2 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFX2 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  ADDFX2 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  ADDFX2 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  ADDFX2 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  ADDFX2 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  ADDFX2 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  ADDFX2 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFX2 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  ADDFX2 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  ADDFX2 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  ADDFX2 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  ADDFX2 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  ADDFX2 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  ADDFX2 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  ADDFX2 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFX2 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  ADDFX2 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  ADDFX2 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  ADDFX2 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  ADDFX2 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  ADDFX2 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  ADDFX2 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  ADDFX2 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  ADDFX2 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFX2 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  ADDFX2 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  ADDFX2 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  ADDFX2 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  ADDFX2 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  ADDFX2 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  ADDFX2 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  ADDFX2 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  ADDFX2 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFX2 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  ADDFX2 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  ADDFX2 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  ADDFX2 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  ADDFX2 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  ADDFX2 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  ADDFX2 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  ADDFX2 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  ADDFX2 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFX2 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  ADDFX2 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  ADDFX2 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  ADDFX2 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  ADDFX2 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  ADDFX2 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  ADDFX2 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  ADDFX2 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  ADDFX2 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  ADDFX2 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  ADDFX2 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  ADDFX2 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  ADDFX2 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  ADDFX2 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  ADDFX2 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  ADDFX2 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  ADDFX2 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  ADDFX2 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  ADDFX2 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFX2 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  ADDFX2 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  ADDFX2 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  ADDFX2 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  ADDFX2 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  ADDFX2 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  ADDFX2 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  ADDFX2 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  ADDFX2 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  ADDFX2 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFX2 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  ADDFX2 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  ADDFX2 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  ADDFX2 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  ADDFX2 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  ADDFX2 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  ADDFX2 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  ADDFX2 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  ADDFX2 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  ADDFX2 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFX2 S2_2_5 ( .A(ab_2__5_), .B(n10), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFX2 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(PRODUCT[11]) );
  ADDFX2 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(PRODUCT[12]) );
  ADDFX2 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT[10]) );
  ADDFX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT[9]) );
  ADDFX2 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT[8]) );
  ADDFX2 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT[7]) );
  ADDFX2 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT[6]) );
  ADDFX2 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT[5]) );
  ADDFX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFX2 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFX2 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFX2 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFX2 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(PRODUCT[15]) );
  ADDFX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFX2 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFX2 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFX2 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFX2 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFX2 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(PRODUCT[14]) );
  ADDFX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFX2 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFX2 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFX2 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFX2 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFX2 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(PRODUCT[13]) );
  ADDFX2 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFX2 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFX2 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFX2 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFX2 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFX2 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFX2 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFX2 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFX2 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFX2 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFX2 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFX2 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFX2 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFX2 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFX2 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFX2 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFX2 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFX2 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFX2 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFX2 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFX2 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFX2 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFX2 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFX2 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFX2 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFX2 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFX2 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFX2 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFX2 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFX2 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFX2 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFX2 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFX2 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFX2 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFX2 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFX2 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFX2 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFX2 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFX2 S2_2_4 ( .A(ab_2__4_), .B(n9), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFX2 S2_2_3 ( .A(ab_2__3_), .B(n13), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFX2 S2_2_2 ( .A(A[2]), .B(n12), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  ADDFX2 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(SUMB_1__1_), .CO(CARRYB_2__0_), 
        .S(PRODUCT[2]) );
  ADDFX2 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFX2 S2_4_4 ( .A(n55), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFX2 S2_3_3 ( .A(n50), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFX2 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT[4]) );
  ADDFX2 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT[3]) );
  ADDFX2 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFX2 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFX2 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFX2 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  ADDFX2 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  AND2X2 U2 ( .A(ab_0__2_), .B(n40), .Y(n7) );
  AND2X2 U3 ( .A(ab_0__1_), .B(ab_1__0_), .Y(n8) );
  AND2X2 U4 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n9) );
  AND2X2 U5 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n10) );
  AND2X2 U6 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n11) );
  AND2X2 U7 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n12) );
  AND2X2 U8 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n13) );
  AND2X2 U9 ( .A(ab_0__8_), .B(ab_1__7_), .Y(n14) );
  AND2X2 U10 ( .A(ab_0__10_), .B(ab_1__9_), .Y(n15) );
  AND2X2 U11 ( .A(ab_0__11_), .B(ab_1__10_), .Y(n16) );
  AND2X2 U12 ( .A(ab_0__12_), .B(ab_1__11_), .Y(n17) );
  AND2X2 U13 ( .A(ab_0__9_), .B(ab_1__8_), .Y(n18) );
  AND2X2 U14 ( .A(ab_0__16_), .B(ab_1__15_), .Y(n19) );
  AND2X2 U15 ( .A(ab_0__13_), .B(ab_1__12_), .Y(n20) );
  AND2X2 U16 ( .A(ab_0__14_), .B(ab_1__13_), .Y(n21) );
  AND2X2 U17 ( .A(ab_0__15_), .B(ab_1__14_), .Y(n22) );
  AND2X2 U18 ( .A(ab_0__17_), .B(ab_1__16_), .Y(n23) );
  AND2X2 U19 ( .A(ab_0__18_), .B(ab_1__17_), .Y(n24) );
  AND2X2 U20 ( .A(ab_0__19_), .B(ab_1__18_), .Y(n25) );
  AND2X2 U21 ( .A(ab_0__20_), .B(ab_1__19_), .Y(n26) );
  AND2X2 U22 ( .A(ab_0__21_), .B(ab_1__20_), .Y(n27) );
  AND2X2 U23 ( .A(ab_0__22_), .B(ab_1__21_), .Y(n28) );
  AND2X2 U24 ( .A(ab_0__23_), .B(ab_1__22_), .Y(n29) );
  AND2X2 U25 ( .A(ab_0__24_), .B(ab_1__23_), .Y(n30) );
  AND2X2 U26 ( .A(ab_0__25_), .B(ab_1__24_), .Y(n31) );
  AND2X2 U27 ( .A(ab_0__26_), .B(ab_1__25_), .Y(n32) );
  AND2X2 U28 ( .A(ab_0__27_), .B(ab_1__26_), .Y(n33) );
  AND2X2 U29 ( .A(ab_0__28_), .B(ab_1__27_), .Y(n34) );
  AND2X2 U30 ( .A(ab_0__29_), .B(ab_1__28_), .Y(n35) );
  AND2X2 U31 ( .A(ab_0__30_), .B(ab_1__29_), .Y(n36) );
  XOR2X1 U32 ( .A(ab_1__0_), .B(ab_0__1_), .Y(PRODUCT[1]) );
  XOR2X1 U33 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X1 U34 ( .A(n40), .B(ab_0__2_), .Y(SUMB_1__1_) );
  XOR2X1 U35 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR2X1 U36 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  XOR2X1 U37 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  INVX1 U38 ( .A(A[2]), .Y(n46) );
  INVX1 U39 ( .A(n50), .Y(n51) );
  INVX1 U40 ( .A(n55), .Y(n57) );
  INVX1 U41 ( .A(A[3]), .Y(n53) );
  INVX1 U42 ( .A(B[2]), .Y(n48) );
  INVX1 U43 ( .A(A[3]), .Y(n54) );
  INVX1 U44 ( .A(n41), .Y(n45) );
  INVX1 U45 ( .A(B[2]), .Y(n47) );
  INVX1 U46 ( .A(n50), .Y(n52) );
  INVX1 U47 ( .A(A[0]), .Y(n39) );
  INVX1 U48 ( .A(A[0]), .Y(n38) );
  INVX1 U49 ( .A(n55), .Y(n58) );
  INVX1 U50 ( .A(n41), .Y(n44) );
  INVX1 U51 ( .A(n40), .Y(n43) );
  INVX1 U52 ( .A(B[2]), .Y(n49) );
  INVX1 U53 ( .A(A[4]), .Y(n59) );
  XOR2X1 U54 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  INVX1 U55 ( .A(n53), .Y(n50) );
  INVX1 U56 ( .A(n56), .Y(n55) );
  INVX1 U57 ( .A(n38), .Y(PRODUCT[0]) );
  XOR2X1 U58 ( .A(ab_1__16_), .B(ab_0__17_), .Y(SUMB_1__16_) );
  XOR2X1 U59 ( .A(ab_1__7_), .B(ab_0__8_), .Y(SUMB_1__7_) );
  XOR2X1 U60 ( .A(ab_1__8_), .B(ab_0__9_), .Y(SUMB_1__8_) );
  XOR2X1 U61 ( .A(ab_1__9_), .B(ab_0__10_), .Y(SUMB_1__9_) );
  XOR2X1 U62 ( .A(ab_1__10_), .B(ab_0__11_), .Y(SUMB_1__10_) );
  XOR2X1 U63 ( .A(ab_1__11_), .B(ab_0__12_), .Y(SUMB_1__11_) );
  XOR2X1 U64 ( .A(ab_1__12_), .B(ab_0__13_), .Y(SUMB_1__12_) );
  XOR2X1 U65 ( .A(ab_1__13_), .B(ab_0__14_), .Y(SUMB_1__13_) );
  XOR2X1 U66 ( .A(ab_1__14_), .B(ab_0__15_), .Y(SUMB_1__14_) );
  XOR2X1 U67 ( .A(ab_1__15_), .B(ab_0__16_), .Y(SUMB_1__15_) );
  INVX1 U68 ( .A(n42), .Y(n40) );
  INVX1 U69 ( .A(n42), .Y(n41) );
  XOR2X1 U70 ( .A(CARRYB_30__0_), .B(SUMB_30__1_), .Y(PRODUCT[31]) );
  INVX1 U71 ( .A(B[1]), .Y(n42) );
  INVX1 U72 ( .A(B[4]), .Y(n56) );
  XOR2X1 U73 ( .A(ab_1__17_), .B(ab_0__18_), .Y(SUMB_1__17_) );
  XOR2X1 U74 ( .A(ab_1__18_), .B(ab_0__19_), .Y(SUMB_1__18_) );
  XOR2X1 U75 ( .A(ab_1__19_), .B(ab_0__20_), .Y(SUMB_1__19_) );
  XOR2X1 U76 ( .A(ab_1__20_), .B(ab_0__21_), .Y(SUMB_1__20_) );
  XOR2X1 U77 ( .A(ab_1__21_), .B(ab_0__22_), .Y(SUMB_1__21_) );
  XOR2X1 U78 ( .A(ab_1__22_), .B(ab_0__23_), .Y(SUMB_1__22_) );
  XOR2X1 U79 ( .A(ab_1__23_), .B(ab_0__24_), .Y(SUMB_1__23_) );
  XOR2X1 U80 ( .A(ab_1__24_), .B(ab_0__25_), .Y(SUMB_1__24_) );
  XOR2X1 U81 ( .A(ab_1__25_), .B(ab_0__26_), .Y(SUMB_1__25_) );
  XOR2X1 U82 ( .A(ab_1__26_), .B(ab_0__27_), .Y(SUMB_1__26_) );
  XOR2X1 U83 ( .A(ab_1__27_), .B(ab_0__28_), .Y(SUMB_1__27_) );
  XOR2X1 U84 ( .A(ab_1__28_), .B(ab_0__29_), .Y(SUMB_1__28_) );
  XOR2X1 U85 ( .A(ab_1__29_), .B(ab_0__30_), .Y(SUMB_1__29_) );
  INVX1 U86 ( .A(B[8]), .Y(n65) );
  INVX1 U87 ( .A(B[12]), .Y(n71) );
  INVX1 U88 ( .A(B[5]), .Y(n60) );
  INVX1 U89 ( .A(B[6]), .Y(n61) );
  INVX1 U90 ( .A(B[7]), .Y(n63) );
  INVX1 U91 ( .A(B[8]), .Y(n64) );
  INVX1 U92 ( .A(B[9]), .Y(n66) );
  INVX1 U93 ( .A(B[10]), .Y(n68) );
  INVX1 U94 ( .A(B[11]), .Y(n70) );
  INVX1 U95 ( .A(B[6]), .Y(n62) );
  INVX1 U96 ( .A(B[13]), .Y(n72) );
  INVX1 U97 ( .A(B[15]), .Y(n74) );
  INVX1 U98 ( .A(B[14]), .Y(n73) );
  INVX1 U99 ( .A(B[9]), .Y(n67) );
  INVX1 U100 ( .A(B[10]), .Y(n69) );
  INVX1 U101 ( .A(B[16]), .Y(n76) );
  INVX1 U102 ( .A(B[17]), .Y(n77) );
  INVX1 U103 ( .A(B[18]), .Y(n78) );
  INVX1 U104 ( .A(B[19]), .Y(n79) );
  INVX1 U105 ( .A(B[20]), .Y(n80) );
  INVX1 U106 ( .A(B[21]), .Y(n81) );
  INVX1 U107 ( .A(B[22]), .Y(n82) );
  INVX1 U108 ( .A(B[23]), .Y(n83) );
  INVX1 U109 ( .A(B[24]), .Y(n84) );
  INVX1 U110 ( .A(B[25]), .Y(n85) );
  INVX1 U111 ( .A(B[26]), .Y(n86) );
  INVX1 U112 ( .A(B[27]), .Y(n87) );
  INVX1 U113 ( .A(B[28]), .Y(n88) );
  INVX1 U114 ( .A(B[29]), .Y(n89) );
  INVX1 U115 ( .A(B[30]), .Y(n75) );
  NOR2X1 U116 ( .A(n66), .B(n65), .Y(ab_9__8_) );
  NOR2X1 U117 ( .A(n67), .B(n63), .Y(ab_9__7_) );
  NOR2X1 U118 ( .A(n66), .B(n62), .Y(ab_9__6_) );
  NOR2X1 U119 ( .A(n66), .B(n60), .Y(ab_9__5_) );
  NOR2X1 U120 ( .A(n66), .B(n59), .Y(ab_9__4_) );
  NOR2X1 U121 ( .A(n66), .B(n53), .Y(ab_9__3_) );
  NOR2X1 U122 ( .A(n66), .B(n47), .Y(ab_9__2_) );
  NOR2X1 U123 ( .A(n67), .B(n82), .Y(ab_9__22_) );
  NOR2X1 U124 ( .A(n67), .B(n81), .Y(ab_9__21_) );
  NOR2X1 U125 ( .A(n66), .B(n80), .Y(ab_9__20_) );
  NOR2X1 U126 ( .A(n66), .B(n45), .Y(ab_9__1_) );
  NOR2X1 U127 ( .A(n67), .B(n79), .Y(ab_9__19_) );
  NOR2X1 U128 ( .A(n66), .B(n78), .Y(ab_9__18_) );
  NOR2X1 U129 ( .A(n67), .B(n77), .Y(ab_9__17_) );
  NOR2X1 U130 ( .A(n67), .B(n76), .Y(ab_9__16_) );
  NOR2X1 U131 ( .A(n66), .B(n74), .Y(ab_9__15_) );
  NOR2X1 U132 ( .A(n67), .B(n73), .Y(ab_9__14_) );
  NOR2X1 U133 ( .A(n66), .B(n72), .Y(ab_9__13_) );
  NOR2X1 U134 ( .A(n67), .B(n71), .Y(ab_9__12_) );
  NOR2X1 U135 ( .A(n66), .B(n70), .Y(ab_9__11_) );
  NOR2X1 U136 ( .A(n67), .B(n69), .Y(ab_9__10_) );
  NOR2X1 U137 ( .A(n66), .B(n39), .Y(ab_9__0_) );
  NOR2X1 U138 ( .A(n66), .B(n65), .Y(ab_8__9_) );
  NOR2X1 U139 ( .A(n63), .B(n65), .Y(ab_8__7_) );
  NOR2X1 U140 ( .A(n62), .B(n65), .Y(ab_8__6_) );
  NOR2X1 U141 ( .A(n60), .B(n65), .Y(ab_8__5_) );
  NOR2X1 U142 ( .A(n59), .B(n65), .Y(ab_8__4_) );
  NOR2X1 U143 ( .A(n53), .B(n65), .Y(ab_8__3_) );
  NOR2X1 U144 ( .A(n47), .B(n65), .Y(ab_8__2_) );
  NOR2X1 U145 ( .A(n83), .B(n65), .Y(ab_8__23_) );
  NOR2X1 U146 ( .A(n82), .B(n65), .Y(ab_8__22_) );
  NOR2X1 U147 ( .A(n81), .B(n65), .Y(ab_8__21_) );
  NOR2X1 U148 ( .A(n80), .B(n65), .Y(ab_8__20_) );
  NOR2X1 U149 ( .A(n45), .B(n65), .Y(ab_8__1_) );
  NOR2X1 U150 ( .A(n79), .B(n65), .Y(ab_8__19_) );
  NOR2X1 U151 ( .A(n78), .B(n65), .Y(ab_8__18_) );
  NOR2X1 U152 ( .A(n77), .B(n65), .Y(ab_8__17_) );
  NOR2X1 U153 ( .A(n76), .B(n65), .Y(ab_8__16_) );
  NOR2X1 U154 ( .A(n74), .B(n65), .Y(ab_8__15_) );
  NOR2X1 U155 ( .A(n73), .B(n65), .Y(ab_8__14_) );
  NOR2X1 U156 ( .A(n72), .B(n65), .Y(ab_8__13_) );
  NOR2X1 U157 ( .A(n71), .B(n65), .Y(ab_8__12_) );
  NOR2X1 U158 ( .A(n70), .B(n65), .Y(ab_8__11_) );
  NOR2X1 U159 ( .A(n69), .B(n65), .Y(ab_8__10_) );
  NOR2X1 U160 ( .A(n39), .B(n65), .Y(ab_8__0_) );
  NOR2X1 U161 ( .A(n66), .B(n63), .Y(ab_7__9_) );
  NOR2X1 U162 ( .A(n65), .B(n63), .Y(ab_7__8_) );
  NOR2X1 U163 ( .A(n62), .B(n63), .Y(ab_7__6_) );
  NOR2X1 U164 ( .A(n60), .B(n63), .Y(ab_7__5_) );
  NOR2X1 U165 ( .A(n59), .B(n63), .Y(ab_7__4_) );
  NOR2X1 U166 ( .A(n53), .B(n63), .Y(ab_7__3_) );
  NOR2X1 U167 ( .A(n47), .B(n63), .Y(ab_7__2_) );
  NOR2X1 U168 ( .A(n84), .B(n63), .Y(ab_7__24_) );
  NOR2X1 U169 ( .A(n83), .B(n63), .Y(ab_7__23_) );
  NOR2X1 U170 ( .A(n82), .B(n63), .Y(ab_7__22_) );
  NOR2X1 U171 ( .A(n81), .B(n63), .Y(ab_7__21_) );
  NOR2X1 U172 ( .A(n80), .B(n63), .Y(ab_7__20_) );
  NOR2X1 U173 ( .A(n45), .B(n63), .Y(ab_7__1_) );
  NOR2X1 U174 ( .A(n79), .B(n63), .Y(ab_7__19_) );
  NOR2X1 U175 ( .A(n78), .B(n63), .Y(ab_7__18_) );
  NOR2X1 U176 ( .A(n77), .B(n63), .Y(ab_7__17_) );
  NOR2X1 U177 ( .A(n76), .B(n63), .Y(ab_7__16_) );
  NOR2X1 U178 ( .A(n74), .B(n63), .Y(ab_7__15_) );
  NOR2X1 U179 ( .A(n73), .B(n63), .Y(ab_7__14_) );
  NOR2X1 U180 ( .A(n72), .B(n63), .Y(ab_7__13_) );
  NOR2X1 U181 ( .A(n71), .B(n63), .Y(ab_7__12_) );
  NOR2X1 U182 ( .A(n70), .B(n63), .Y(ab_7__11_) );
  NOR2X1 U183 ( .A(n69), .B(n63), .Y(ab_7__10_) );
  NOR2X1 U184 ( .A(n39), .B(n63), .Y(ab_7__0_) );
  NOR2X1 U185 ( .A(n66), .B(n62), .Y(ab_6__9_) );
  NOR2X1 U186 ( .A(n65), .B(n62), .Y(ab_6__8_) );
  NOR2X1 U187 ( .A(n63), .B(n62), .Y(ab_6__7_) );
  NOR2X1 U188 ( .A(n60), .B(n62), .Y(ab_6__5_) );
  NOR2X1 U189 ( .A(n58), .B(n62), .Y(ab_6__4_) );
  NOR2X1 U190 ( .A(n53), .B(n62), .Y(ab_6__3_) );
  NOR2X1 U191 ( .A(n47), .B(n62), .Y(ab_6__2_) );
  NOR2X1 U192 ( .A(n85), .B(n62), .Y(ab_6__25_) );
  NOR2X1 U193 ( .A(n84), .B(n62), .Y(ab_6__24_) );
  NOR2X1 U194 ( .A(n83), .B(n62), .Y(ab_6__23_) );
  NOR2X1 U195 ( .A(n82), .B(n62), .Y(ab_6__22_) );
  NOR2X1 U196 ( .A(n81), .B(n62), .Y(ab_6__21_) );
  NOR2X1 U197 ( .A(n80), .B(n62), .Y(ab_6__20_) );
  NOR2X1 U198 ( .A(n45), .B(n62), .Y(ab_6__1_) );
  NOR2X1 U199 ( .A(n79), .B(n62), .Y(ab_6__19_) );
  NOR2X1 U200 ( .A(n78), .B(n62), .Y(ab_6__18_) );
  NOR2X1 U201 ( .A(n77), .B(n62), .Y(ab_6__17_) );
  NOR2X1 U202 ( .A(n76), .B(n62), .Y(ab_6__16_) );
  NOR2X1 U203 ( .A(n74), .B(n62), .Y(ab_6__15_) );
  NOR2X1 U204 ( .A(n73), .B(n62), .Y(ab_6__14_) );
  NOR2X1 U205 ( .A(n72), .B(n62), .Y(ab_6__13_) );
  NOR2X1 U206 ( .A(n71), .B(n62), .Y(ab_6__12_) );
  NOR2X1 U207 ( .A(n70), .B(n62), .Y(ab_6__11_) );
  NOR2X1 U208 ( .A(n69), .B(n62), .Y(ab_6__10_) );
  NOR2X1 U209 ( .A(n39), .B(n62), .Y(ab_6__0_) );
  NOR2X1 U210 ( .A(n66), .B(n60), .Y(ab_5__9_) );
  NOR2X1 U211 ( .A(n65), .B(n60), .Y(ab_5__8_) );
  NOR2X1 U212 ( .A(n63), .B(n60), .Y(ab_5__7_) );
  NOR2X1 U213 ( .A(n62), .B(n60), .Y(ab_5__6_) );
  NOR2X1 U214 ( .A(n58), .B(n60), .Y(ab_5__4_) );
  NOR2X1 U215 ( .A(n52), .B(n60), .Y(ab_5__3_) );
  NOR2X1 U216 ( .A(n47), .B(n60), .Y(ab_5__2_) );
  NOR2X1 U217 ( .A(n86), .B(n60), .Y(ab_5__26_) );
  NOR2X1 U218 ( .A(n85), .B(n60), .Y(ab_5__25_) );
  NOR2X1 U219 ( .A(n84), .B(n60), .Y(ab_5__24_) );
  NOR2X1 U220 ( .A(n83), .B(n60), .Y(ab_5__23_) );
  NOR2X1 U221 ( .A(n82), .B(n60), .Y(ab_5__22_) );
  NOR2X1 U222 ( .A(n81), .B(n60), .Y(ab_5__21_) );
  NOR2X1 U223 ( .A(n80), .B(n60), .Y(ab_5__20_) );
  NOR2X1 U224 ( .A(n45), .B(n60), .Y(ab_5__1_) );
  NOR2X1 U225 ( .A(n79), .B(n60), .Y(ab_5__19_) );
  NOR2X1 U226 ( .A(n78), .B(n60), .Y(ab_5__18_) );
  NOR2X1 U227 ( .A(n77), .B(n60), .Y(ab_5__17_) );
  NOR2X1 U228 ( .A(n76), .B(n60), .Y(ab_5__16_) );
  NOR2X1 U229 ( .A(n74), .B(n60), .Y(ab_5__15_) );
  NOR2X1 U230 ( .A(n73), .B(n60), .Y(ab_5__14_) );
  NOR2X1 U231 ( .A(n72), .B(n60), .Y(ab_5__13_) );
  NOR2X1 U232 ( .A(n71), .B(n60), .Y(ab_5__12_) );
  NOR2X1 U233 ( .A(n70), .B(n60), .Y(ab_5__11_) );
  NOR2X1 U234 ( .A(n69), .B(n60), .Y(ab_5__10_) );
  NOR2X1 U235 ( .A(n39), .B(n60), .Y(ab_5__0_) );
  NOR2X1 U236 ( .A(n66), .B(n59), .Y(ab_4__9_) );
  NOR2X1 U237 ( .A(n65), .B(n59), .Y(ab_4__8_) );
  NOR2X1 U238 ( .A(n63), .B(n59), .Y(ab_4__7_) );
  NOR2X1 U239 ( .A(n62), .B(n59), .Y(ab_4__6_) );
  NOR2X1 U240 ( .A(n60), .B(n59), .Y(ab_4__5_) );
  NOR2X1 U241 ( .A(n52), .B(n59), .Y(ab_4__3_) );
  NOR2X1 U242 ( .A(n49), .B(n59), .Y(ab_4__2_) );
  NOR2X1 U243 ( .A(n87), .B(n59), .Y(ab_4__27_) );
  NOR2X1 U244 ( .A(n86), .B(n59), .Y(ab_4__26_) );
  NOR2X1 U245 ( .A(n85), .B(n59), .Y(ab_4__25_) );
  NOR2X1 U246 ( .A(n84), .B(n59), .Y(ab_4__24_) );
  NOR2X1 U247 ( .A(n83), .B(n59), .Y(ab_4__23_) );
  NOR2X1 U248 ( .A(n82), .B(n59), .Y(ab_4__22_) );
  NOR2X1 U249 ( .A(n81), .B(n59), .Y(ab_4__21_) );
  NOR2X1 U250 ( .A(n80), .B(n59), .Y(ab_4__20_) );
  NOR2X1 U251 ( .A(n45), .B(n59), .Y(ab_4__1_) );
  NOR2X1 U252 ( .A(n79), .B(n59), .Y(ab_4__19_) );
  NOR2X1 U253 ( .A(n78), .B(n59), .Y(ab_4__18_) );
  NOR2X1 U254 ( .A(n77), .B(n59), .Y(ab_4__17_) );
  NOR2X1 U255 ( .A(n76), .B(n59), .Y(ab_4__16_) );
  NOR2X1 U256 ( .A(n74), .B(n59), .Y(ab_4__15_) );
  NOR2X1 U257 ( .A(n73), .B(n59), .Y(ab_4__14_) );
  NOR2X1 U258 ( .A(n72), .B(n59), .Y(ab_4__13_) );
  NOR2X1 U259 ( .A(n71), .B(n59), .Y(ab_4__12_) );
  NOR2X1 U260 ( .A(n70), .B(n59), .Y(ab_4__11_) );
  NOR2X1 U261 ( .A(n69), .B(n59), .Y(ab_4__10_) );
  NOR2X1 U262 ( .A(n39), .B(n59), .Y(ab_4__0_) );
  NOR2X1 U263 ( .A(n66), .B(n54), .Y(ab_3__9_) );
  NOR2X1 U264 ( .A(n65), .B(n54), .Y(ab_3__8_) );
  NOR2X1 U265 ( .A(n63), .B(n54), .Y(ab_3__7_) );
  NOR2X1 U266 ( .A(n62), .B(n54), .Y(ab_3__6_) );
  NOR2X1 U267 ( .A(n60), .B(n54), .Y(ab_3__5_) );
  NOR2X1 U268 ( .A(n58), .B(n54), .Y(ab_3__4_) );
  NOR2X1 U269 ( .A(n49), .B(n54), .Y(ab_3__2_) );
  NOR2X1 U270 ( .A(n88), .B(n54), .Y(ab_3__28_) );
  NOR2X1 U271 ( .A(n87), .B(n54), .Y(ab_3__27_) );
  NOR2X1 U272 ( .A(n86), .B(n54), .Y(ab_3__26_) );
  NOR2X1 U273 ( .A(n85), .B(n54), .Y(ab_3__25_) );
  NOR2X1 U274 ( .A(n84), .B(n54), .Y(ab_3__24_) );
  NOR2X1 U275 ( .A(n83), .B(n54), .Y(ab_3__23_) );
  NOR2X1 U276 ( .A(n82), .B(n54), .Y(ab_3__22_) );
  NOR2X1 U277 ( .A(n81), .B(n54), .Y(ab_3__21_) );
  NOR2X1 U278 ( .A(n80), .B(n54), .Y(ab_3__20_) );
  NOR2X1 U279 ( .A(n44), .B(n54), .Y(ab_3__1_) );
  NOR2X1 U280 ( .A(n79), .B(n54), .Y(ab_3__19_) );
  NOR2X1 U281 ( .A(n78), .B(n53), .Y(ab_3__18_) );
  NOR2X1 U282 ( .A(n77), .B(n53), .Y(ab_3__17_) );
  NOR2X1 U283 ( .A(n76), .B(n53), .Y(ab_3__16_) );
  NOR2X1 U284 ( .A(n74), .B(n53), .Y(ab_3__15_) );
  NOR2X1 U285 ( .A(n73), .B(n53), .Y(ab_3__14_) );
  NOR2X1 U286 ( .A(n72), .B(n53), .Y(ab_3__13_) );
  NOR2X1 U287 ( .A(n71), .B(n53), .Y(ab_3__12_) );
  NOR2X1 U288 ( .A(n70), .B(n53), .Y(ab_3__11_) );
  NOR2X1 U289 ( .A(n69), .B(n53), .Y(ab_3__10_) );
  NOR2X1 U290 ( .A(n39), .B(n53), .Y(ab_3__0_) );
  NOR2X1 U291 ( .A(n44), .B(n75), .Y(ab_30__1_) );
  NOR2X1 U292 ( .A(n39), .B(n75), .Y(ab_30__0_) );
  NOR2X1 U293 ( .A(n66), .B(n49), .Y(ab_2__9_) );
  NOR2X1 U294 ( .A(n65), .B(n49), .Y(ab_2__8_) );
  NOR2X1 U295 ( .A(n63), .B(n49), .Y(ab_2__7_) );
  NOR2X1 U296 ( .A(n62), .B(n49), .Y(ab_2__6_) );
  NOR2X1 U297 ( .A(n60), .B(n49), .Y(ab_2__5_) );
  NOR2X1 U298 ( .A(n58), .B(n49), .Y(ab_2__4_) );
  NOR2X1 U299 ( .A(n52), .B(n49), .Y(ab_2__3_) );
  NOR2X1 U300 ( .A(n89), .B(n48), .Y(ab_2__29_) );
  NOR2X1 U301 ( .A(n88), .B(n48), .Y(ab_2__28_) );
  NOR2X1 U302 ( .A(n87), .B(n48), .Y(ab_2__27_) );
  NOR2X1 U303 ( .A(n86), .B(n48), .Y(ab_2__26_) );
  NOR2X1 U304 ( .A(n85), .B(n48), .Y(ab_2__25_) );
  NOR2X1 U305 ( .A(n84), .B(n48), .Y(ab_2__24_) );
  NOR2X1 U306 ( .A(n83), .B(n48), .Y(ab_2__23_) );
  NOR2X1 U307 ( .A(n82), .B(n48), .Y(ab_2__22_) );
  NOR2X1 U308 ( .A(n81), .B(n48), .Y(ab_2__21_) );
  NOR2X1 U309 ( .A(n80), .B(n48), .Y(ab_2__20_) );
  NOR2X1 U310 ( .A(n44), .B(n48), .Y(ab_2__1_) );
  NOR2X1 U311 ( .A(n79), .B(n48), .Y(ab_2__19_) );
  NOR2X1 U312 ( .A(n78), .B(n48), .Y(ab_2__18_) );
  NOR2X1 U313 ( .A(n77), .B(n48), .Y(ab_2__17_) );
  NOR2X1 U314 ( .A(n76), .B(n47), .Y(ab_2__16_) );
  NOR2X1 U315 ( .A(n74), .B(n47), .Y(ab_2__15_) );
  NOR2X1 U316 ( .A(n73), .B(n47), .Y(ab_2__14_) );
  NOR2X1 U317 ( .A(n72), .B(n47), .Y(ab_2__13_) );
  NOR2X1 U318 ( .A(n71), .B(n47), .Y(ab_2__12_) );
  NOR2X1 U319 ( .A(n70), .B(n47), .Y(ab_2__11_) );
  NOR2X1 U320 ( .A(n69), .B(n47), .Y(ab_2__10_) );
  NOR2X1 U321 ( .A(n39), .B(n47), .Y(ab_2__0_) );
  NOR2X1 U322 ( .A(n49), .B(n89), .Y(ab_29__2_) );
  NOR2X1 U323 ( .A(n44), .B(n89), .Y(ab_29__1_) );
  NOR2X1 U324 ( .A(n39), .B(n89), .Y(ab_29__0_) );
  NOR2X1 U325 ( .A(n52), .B(n88), .Y(ab_28__3_) );
  NOR2X1 U326 ( .A(n49), .B(n88), .Y(ab_28__2_) );
  NOR2X1 U327 ( .A(n44), .B(n88), .Y(ab_28__1_) );
  NOR2X1 U328 ( .A(n39), .B(n88), .Y(ab_28__0_) );
  NOR2X1 U329 ( .A(n58), .B(n87), .Y(ab_27__4_) );
  NOR2X1 U330 ( .A(n52), .B(n87), .Y(ab_27__3_) );
  NOR2X1 U331 ( .A(n49), .B(n87), .Y(ab_27__2_) );
  NOR2X1 U332 ( .A(n44), .B(n87), .Y(ab_27__1_) );
  NOR2X1 U333 ( .A(n39), .B(n87), .Y(ab_27__0_) );
  NOR2X1 U334 ( .A(n60), .B(n86), .Y(ab_26__5_) );
  NOR2X1 U335 ( .A(n58), .B(n86), .Y(ab_26__4_) );
  NOR2X1 U336 ( .A(n52), .B(n86), .Y(ab_26__3_) );
  NOR2X1 U337 ( .A(n49), .B(n86), .Y(ab_26__2_) );
  NOR2X1 U338 ( .A(n44), .B(n86), .Y(ab_26__1_) );
  NOR2X1 U339 ( .A(n39), .B(n86), .Y(ab_26__0_) );
  NOR2X1 U340 ( .A(n62), .B(n85), .Y(ab_25__6_) );
  NOR2X1 U341 ( .A(n60), .B(n85), .Y(ab_25__5_) );
  NOR2X1 U342 ( .A(n58), .B(n85), .Y(ab_25__4_) );
  NOR2X1 U343 ( .A(n52), .B(n85), .Y(ab_25__3_) );
  NOR2X1 U344 ( .A(n49), .B(n85), .Y(ab_25__2_) );
  NOR2X1 U345 ( .A(n44), .B(n85), .Y(ab_25__1_) );
  NOR2X1 U346 ( .A(n39), .B(n85), .Y(ab_25__0_) );
  NOR2X1 U347 ( .A(n63), .B(n84), .Y(ab_24__7_) );
  NOR2X1 U348 ( .A(n62), .B(n84), .Y(ab_24__6_) );
  NOR2X1 U349 ( .A(n60), .B(n84), .Y(ab_24__5_) );
  NOR2X1 U350 ( .A(n58), .B(n84), .Y(ab_24__4_) );
  NOR2X1 U351 ( .A(n52), .B(n84), .Y(ab_24__3_) );
  NOR2X1 U352 ( .A(n49), .B(n84), .Y(ab_24__2_) );
  NOR2X1 U353 ( .A(n44), .B(n84), .Y(ab_24__1_) );
  NOR2X1 U354 ( .A(n39), .B(n84), .Y(ab_24__0_) );
  NOR2X1 U355 ( .A(n65), .B(n83), .Y(ab_23__8_) );
  NOR2X1 U356 ( .A(n63), .B(n83), .Y(ab_23__7_) );
  NOR2X1 U357 ( .A(n62), .B(n83), .Y(ab_23__6_) );
  NOR2X1 U358 ( .A(n60), .B(n83), .Y(ab_23__5_) );
  NOR2X1 U359 ( .A(n58), .B(n83), .Y(ab_23__4_) );
  NOR2X1 U360 ( .A(n52), .B(n83), .Y(ab_23__3_) );
  NOR2X1 U361 ( .A(n49), .B(n83), .Y(ab_23__2_) );
  NOR2X1 U362 ( .A(n44), .B(n83), .Y(ab_23__1_) );
  NOR2X1 U363 ( .A(n39), .B(n83), .Y(ab_23__0_) );
  NOR2X1 U364 ( .A(n66), .B(n82), .Y(ab_22__9_) );
  NOR2X1 U365 ( .A(n65), .B(n82), .Y(ab_22__8_) );
  NOR2X1 U366 ( .A(n63), .B(n82), .Y(ab_22__7_) );
  NOR2X1 U367 ( .A(n62), .B(n82), .Y(ab_22__6_) );
  NOR2X1 U368 ( .A(n60), .B(n82), .Y(ab_22__5_) );
  NOR2X1 U369 ( .A(n58), .B(n82), .Y(ab_22__4_) );
  NOR2X1 U370 ( .A(n52), .B(n82), .Y(ab_22__3_) );
  NOR2X1 U371 ( .A(n49), .B(n82), .Y(ab_22__2_) );
  NOR2X1 U372 ( .A(n44), .B(n82), .Y(ab_22__1_) );
  NOR2X1 U373 ( .A(n39), .B(n82), .Y(ab_22__0_) );
  NOR2X1 U374 ( .A(n66), .B(n81), .Y(ab_21__9_) );
  NOR2X1 U375 ( .A(n65), .B(n81), .Y(ab_21__8_) );
  NOR2X1 U376 ( .A(n63), .B(n81), .Y(ab_21__7_) );
  NOR2X1 U377 ( .A(n62), .B(n81), .Y(ab_21__6_) );
  NOR2X1 U378 ( .A(n60), .B(n81), .Y(ab_21__5_) );
  NOR2X1 U379 ( .A(n58), .B(n81), .Y(ab_21__4_) );
  NOR2X1 U380 ( .A(n52), .B(n81), .Y(ab_21__3_) );
  NOR2X1 U381 ( .A(n49), .B(n81), .Y(ab_21__2_) );
  NOR2X1 U382 ( .A(n44), .B(n81), .Y(ab_21__1_) );
  NOR2X1 U383 ( .A(n69), .B(n81), .Y(ab_21__10_) );
  NOR2X1 U384 ( .A(n39), .B(n81), .Y(ab_21__0_) );
  NOR2X1 U385 ( .A(n66), .B(n80), .Y(ab_20__9_) );
  NOR2X1 U386 ( .A(n65), .B(n80), .Y(ab_20__8_) );
  NOR2X1 U387 ( .A(n63), .B(n80), .Y(ab_20__7_) );
  NOR2X1 U388 ( .A(n62), .B(n80), .Y(ab_20__6_) );
  NOR2X1 U389 ( .A(n60), .B(n80), .Y(ab_20__5_) );
  NOR2X1 U390 ( .A(n58), .B(n80), .Y(ab_20__4_) );
  NOR2X1 U391 ( .A(n52), .B(n80), .Y(ab_20__3_) );
  NOR2X1 U392 ( .A(n49), .B(n80), .Y(ab_20__2_) );
  NOR2X1 U393 ( .A(n43), .B(n80), .Y(ab_20__1_) );
  NOR2X1 U394 ( .A(n70), .B(n80), .Y(ab_20__11_) );
  NOR2X1 U395 ( .A(n68), .B(n80), .Y(ab_20__10_) );
  NOR2X1 U396 ( .A(n38), .B(n80), .Y(ab_20__0_) );
  NOR2X1 U397 ( .A(n66), .B(n45), .Y(ab_1__9_) );
  NOR2X1 U398 ( .A(n64), .B(n44), .Y(ab_1__8_) );
  NOR2X1 U399 ( .A(n63), .B(n44), .Y(ab_1__7_) );
  NOR2X1 U400 ( .A(n61), .B(n44), .Y(ab_1__6_) );
  NOR2X1 U401 ( .A(n60), .B(n44), .Y(ab_1__5_) );
  NOR2X1 U402 ( .A(n57), .B(n44), .Y(ab_1__4_) );
  NOR2X1 U403 ( .A(n51), .B(n44), .Y(ab_1__3_) );
  NOR2X1 U404 ( .A(n75), .B(n44), .Y(ab_1__30_) );
  NOR2X1 U405 ( .A(n46), .B(n44), .Y(ab_1__2_) );
  NOR2X1 U406 ( .A(n89), .B(n44), .Y(ab_1__29_) );
  NOR2X1 U407 ( .A(n88), .B(n45), .Y(ab_1__28_) );
  NOR2X1 U408 ( .A(n87), .B(n44), .Y(ab_1__27_) );
  NOR2X1 U409 ( .A(n86), .B(n43), .Y(ab_1__26_) );
  NOR2X1 U410 ( .A(n85), .B(n44), .Y(ab_1__25_) );
  NOR2X1 U411 ( .A(n84), .B(n44), .Y(ab_1__24_) );
  NOR2X1 U412 ( .A(n83), .B(n45), .Y(ab_1__23_) );
  NOR2X1 U413 ( .A(n82), .B(n44), .Y(ab_1__22_) );
  NOR2X1 U414 ( .A(n81), .B(n44), .Y(ab_1__21_) );
  NOR2X1 U415 ( .A(n80), .B(n44), .Y(ab_1__20_) );
  NOR2X1 U416 ( .A(n79), .B(n45), .Y(ab_1__19_) );
  NOR2X1 U417 ( .A(n78), .B(n44), .Y(ab_1__18_) );
  NOR2X1 U418 ( .A(n77), .B(n45), .Y(ab_1__17_) );
  NOR2X1 U419 ( .A(n76), .B(n44), .Y(ab_1__16_) );
  NOR2X1 U420 ( .A(n74), .B(n45), .Y(ab_1__15_) );
  NOR2X1 U421 ( .A(n73), .B(n45), .Y(ab_1__14_) );
  NOR2X1 U422 ( .A(n72), .B(n45), .Y(ab_1__13_) );
  NOR2X1 U423 ( .A(n71), .B(n45), .Y(ab_1__12_) );
  NOR2X1 U424 ( .A(n70), .B(n45), .Y(ab_1__11_) );
  NOR2X1 U425 ( .A(n68), .B(n45), .Y(ab_1__10_) );
  NOR2X1 U426 ( .A(n38), .B(n45), .Y(ab_1__0_) );
  NOR2X1 U427 ( .A(n66), .B(n79), .Y(ab_19__9_) );
  NOR2X1 U428 ( .A(n64), .B(n79), .Y(ab_19__8_) );
  NOR2X1 U429 ( .A(n63), .B(n79), .Y(ab_19__7_) );
  NOR2X1 U430 ( .A(n61), .B(n79), .Y(ab_19__6_) );
  NOR2X1 U431 ( .A(n60), .B(n79), .Y(ab_19__5_) );
  NOR2X1 U432 ( .A(n57), .B(n79), .Y(ab_19__4_) );
  NOR2X1 U433 ( .A(n51), .B(n79), .Y(ab_19__3_) );
  NOR2X1 U434 ( .A(n46), .B(n79), .Y(ab_19__2_) );
  NOR2X1 U435 ( .A(n43), .B(n79), .Y(ab_19__1_) );
  NOR2X1 U436 ( .A(n71), .B(n79), .Y(ab_19__12_) );
  NOR2X1 U437 ( .A(n70), .B(n79), .Y(ab_19__11_) );
  NOR2X1 U438 ( .A(n68), .B(n79), .Y(ab_19__10_) );
  NOR2X1 U439 ( .A(n38), .B(n79), .Y(ab_19__0_) );
  NOR2X1 U440 ( .A(n66), .B(n78), .Y(ab_18__9_) );
  NOR2X1 U441 ( .A(n64), .B(n78), .Y(ab_18__8_) );
  NOR2X1 U442 ( .A(n63), .B(n78), .Y(ab_18__7_) );
  NOR2X1 U443 ( .A(n61), .B(n78), .Y(ab_18__6_) );
  NOR2X1 U444 ( .A(n60), .B(n78), .Y(ab_18__5_) );
  NOR2X1 U445 ( .A(n57), .B(n78), .Y(ab_18__4_) );
  NOR2X1 U446 ( .A(n51), .B(n78), .Y(ab_18__3_) );
  NOR2X1 U447 ( .A(n46), .B(n78), .Y(ab_18__2_) );
  NOR2X1 U448 ( .A(n43), .B(n78), .Y(ab_18__1_) );
  NOR2X1 U449 ( .A(n72), .B(n78), .Y(ab_18__13_) );
  NOR2X1 U450 ( .A(n71), .B(n78), .Y(ab_18__12_) );
  NOR2X1 U451 ( .A(n70), .B(n78), .Y(ab_18__11_) );
  NOR2X1 U452 ( .A(n68), .B(n78), .Y(ab_18__10_) );
  NOR2X1 U453 ( .A(n38), .B(n78), .Y(ab_18__0_) );
  NOR2X1 U454 ( .A(n66), .B(n77), .Y(ab_17__9_) );
  NOR2X1 U455 ( .A(n64), .B(n77), .Y(ab_17__8_) );
  NOR2X1 U456 ( .A(n63), .B(n77), .Y(ab_17__7_) );
  NOR2X1 U457 ( .A(n61), .B(n77), .Y(ab_17__6_) );
  NOR2X1 U458 ( .A(n60), .B(n77), .Y(ab_17__5_) );
  NOR2X1 U459 ( .A(n57), .B(n77), .Y(ab_17__4_) );
  NOR2X1 U460 ( .A(n51), .B(n77), .Y(ab_17__3_) );
  NOR2X1 U461 ( .A(n46), .B(n77), .Y(ab_17__2_) );
  NOR2X1 U462 ( .A(n43), .B(n77), .Y(ab_17__1_) );
  NOR2X1 U463 ( .A(n73), .B(n77), .Y(ab_17__14_) );
  NOR2X1 U464 ( .A(n72), .B(n77), .Y(ab_17__13_) );
  NOR2X1 U465 ( .A(n71), .B(n77), .Y(ab_17__12_) );
  NOR2X1 U466 ( .A(n70), .B(n77), .Y(ab_17__11_) );
  NOR2X1 U467 ( .A(n68), .B(n77), .Y(ab_17__10_) );
  NOR2X1 U468 ( .A(n38), .B(n77), .Y(ab_17__0_) );
  NOR2X1 U469 ( .A(n67), .B(n76), .Y(ab_16__9_) );
  NOR2X1 U470 ( .A(n64), .B(n76), .Y(ab_16__8_) );
  NOR2X1 U471 ( .A(n63), .B(n76), .Y(ab_16__7_) );
  NOR2X1 U472 ( .A(n61), .B(n76), .Y(ab_16__6_) );
  NOR2X1 U473 ( .A(n60), .B(n76), .Y(ab_16__5_) );
  NOR2X1 U474 ( .A(n57), .B(n76), .Y(ab_16__4_) );
  NOR2X1 U475 ( .A(n51), .B(n76), .Y(ab_16__3_) );
  NOR2X1 U476 ( .A(n46), .B(n76), .Y(ab_16__2_) );
  NOR2X1 U477 ( .A(n43), .B(n76), .Y(ab_16__1_) );
  NOR2X1 U478 ( .A(n74), .B(n76), .Y(ab_16__15_) );
  NOR2X1 U479 ( .A(n73), .B(n76), .Y(ab_16__14_) );
  NOR2X1 U480 ( .A(n72), .B(n76), .Y(ab_16__13_) );
  NOR2X1 U481 ( .A(n71), .B(n76), .Y(ab_16__12_) );
  NOR2X1 U482 ( .A(n70), .B(n76), .Y(ab_16__11_) );
  NOR2X1 U483 ( .A(n68), .B(n76), .Y(ab_16__10_) );
  NOR2X1 U484 ( .A(n38), .B(n76), .Y(ab_16__0_) );
  NOR2X1 U485 ( .A(n67), .B(n74), .Y(ab_15__9_) );
  NOR2X1 U486 ( .A(n64), .B(n74), .Y(ab_15__8_) );
  NOR2X1 U487 ( .A(n63), .B(n74), .Y(ab_15__7_) );
  NOR2X1 U488 ( .A(n61), .B(n74), .Y(ab_15__6_) );
  NOR2X1 U489 ( .A(n60), .B(n74), .Y(ab_15__5_) );
  NOR2X1 U490 ( .A(n57), .B(n74), .Y(ab_15__4_) );
  NOR2X1 U491 ( .A(n51), .B(n74), .Y(ab_15__3_) );
  NOR2X1 U492 ( .A(n46), .B(n74), .Y(ab_15__2_) );
  NOR2X1 U493 ( .A(n43), .B(n74), .Y(ab_15__1_) );
  NOR2X1 U494 ( .A(n76), .B(n74), .Y(ab_15__16_) );
  NOR2X1 U495 ( .A(n73), .B(n74), .Y(ab_15__14_) );
  NOR2X1 U496 ( .A(n72), .B(n74), .Y(ab_15__13_) );
  NOR2X1 U497 ( .A(n71), .B(n74), .Y(ab_15__12_) );
  NOR2X1 U498 ( .A(n70), .B(n74), .Y(ab_15__11_) );
  NOR2X1 U499 ( .A(n68), .B(n74), .Y(ab_15__10_) );
  NOR2X1 U500 ( .A(n38), .B(n74), .Y(ab_15__0_) );
  NOR2X1 U501 ( .A(n67), .B(n73), .Y(ab_14__9_) );
  NOR2X1 U502 ( .A(n64), .B(n73), .Y(ab_14__8_) );
  NOR2X1 U503 ( .A(n63), .B(n73), .Y(ab_14__7_) );
  NOR2X1 U504 ( .A(n61), .B(n73), .Y(ab_14__6_) );
  NOR2X1 U505 ( .A(n60), .B(n73), .Y(ab_14__5_) );
  NOR2X1 U506 ( .A(n57), .B(n73), .Y(ab_14__4_) );
  NOR2X1 U507 ( .A(n51), .B(n73), .Y(ab_14__3_) );
  NOR2X1 U508 ( .A(n46), .B(n73), .Y(ab_14__2_) );
  NOR2X1 U509 ( .A(n43), .B(n73), .Y(ab_14__1_) );
  NOR2X1 U510 ( .A(n77), .B(n73), .Y(ab_14__17_) );
  NOR2X1 U511 ( .A(n76), .B(n73), .Y(ab_14__16_) );
  NOR2X1 U512 ( .A(n74), .B(n73), .Y(ab_14__15_) );
  NOR2X1 U513 ( .A(n72), .B(n73), .Y(ab_14__13_) );
  NOR2X1 U514 ( .A(n71), .B(n73), .Y(ab_14__12_) );
  NOR2X1 U515 ( .A(n70), .B(n73), .Y(ab_14__11_) );
  NOR2X1 U516 ( .A(n68), .B(n73), .Y(ab_14__10_) );
  NOR2X1 U517 ( .A(n38), .B(n73), .Y(ab_14__0_) );
  NOR2X1 U518 ( .A(n67), .B(n72), .Y(ab_13__9_) );
  NOR2X1 U519 ( .A(n64), .B(n72), .Y(ab_13__8_) );
  NOR2X1 U520 ( .A(n63), .B(n72), .Y(ab_13__7_) );
  NOR2X1 U521 ( .A(n61), .B(n72), .Y(ab_13__6_) );
  NOR2X1 U522 ( .A(n60), .B(n72), .Y(ab_13__5_) );
  NOR2X1 U523 ( .A(n57), .B(n72), .Y(ab_13__4_) );
  NOR2X1 U524 ( .A(n51), .B(n72), .Y(ab_13__3_) );
  NOR2X1 U525 ( .A(n46), .B(n72), .Y(ab_13__2_) );
  NOR2X1 U526 ( .A(n43), .B(n72), .Y(ab_13__1_) );
  NOR2X1 U527 ( .A(n78), .B(n72), .Y(ab_13__18_) );
  NOR2X1 U528 ( .A(n77), .B(n72), .Y(ab_13__17_) );
  NOR2X1 U529 ( .A(n76), .B(n72), .Y(ab_13__16_) );
  NOR2X1 U530 ( .A(n74), .B(n72), .Y(ab_13__15_) );
  NOR2X1 U531 ( .A(n73), .B(n72), .Y(ab_13__14_) );
  NOR2X1 U532 ( .A(n71), .B(n72), .Y(ab_13__12_) );
  NOR2X1 U533 ( .A(n70), .B(n72), .Y(ab_13__11_) );
  NOR2X1 U534 ( .A(n68), .B(n72), .Y(ab_13__10_) );
  NOR2X1 U535 ( .A(n38), .B(n72), .Y(ab_13__0_) );
  NOR2X1 U536 ( .A(n67), .B(n71), .Y(ab_12__9_) );
  NOR2X1 U537 ( .A(n64), .B(n71), .Y(ab_12__8_) );
  NOR2X1 U538 ( .A(n63), .B(n71), .Y(ab_12__7_) );
  NOR2X1 U539 ( .A(n61), .B(n71), .Y(ab_12__6_) );
  NOR2X1 U540 ( .A(n60), .B(n71), .Y(ab_12__5_) );
  NOR2X1 U541 ( .A(n57), .B(n71), .Y(ab_12__4_) );
  NOR2X1 U542 ( .A(n51), .B(n71), .Y(ab_12__3_) );
  NOR2X1 U543 ( .A(n46), .B(n71), .Y(ab_12__2_) );
  NOR2X1 U544 ( .A(n43), .B(n71), .Y(ab_12__1_) );
  NOR2X1 U545 ( .A(n79), .B(n71), .Y(ab_12__19_) );
  NOR2X1 U546 ( .A(n78), .B(n71), .Y(ab_12__18_) );
  NOR2X1 U547 ( .A(n77), .B(n71), .Y(ab_12__17_) );
  NOR2X1 U548 ( .A(n76), .B(n71), .Y(ab_12__16_) );
  NOR2X1 U549 ( .A(n74), .B(n71), .Y(ab_12__15_) );
  NOR2X1 U550 ( .A(n73), .B(n71), .Y(ab_12__14_) );
  NOR2X1 U551 ( .A(n72), .B(n71), .Y(ab_12__13_) );
  NOR2X1 U552 ( .A(n70), .B(n71), .Y(ab_12__11_) );
  NOR2X1 U553 ( .A(n68), .B(n71), .Y(ab_12__10_) );
  NOR2X1 U554 ( .A(n38), .B(n71), .Y(ab_12__0_) );
  NOR2X1 U555 ( .A(n67), .B(n70), .Y(ab_11__9_) );
  NOR2X1 U556 ( .A(n64), .B(n70), .Y(ab_11__8_) );
  NOR2X1 U557 ( .A(n63), .B(n70), .Y(ab_11__7_) );
  NOR2X1 U558 ( .A(n61), .B(n70), .Y(ab_11__6_) );
  NOR2X1 U559 ( .A(n60), .B(n70), .Y(ab_11__5_) );
  NOR2X1 U560 ( .A(n57), .B(n70), .Y(ab_11__4_) );
  NOR2X1 U561 ( .A(n51), .B(n70), .Y(ab_11__3_) );
  NOR2X1 U562 ( .A(n46), .B(n70), .Y(ab_11__2_) );
  NOR2X1 U563 ( .A(n80), .B(n70), .Y(ab_11__20_) );
  NOR2X1 U564 ( .A(n43), .B(n70), .Y(ab_11__1_) );
  NOR2X1 U565 ( .A(n79), .B(n70), .Y(ab_11__19_) );
  NOR2X1 U566 ( .A(n78), .B(n70), .Y(ab_11__18_) );
  NOR2X1 U567 ( .A(n77), .B(n70), .Y(ab_11__17_) );
  NOR2X1 U568 ( .A(n76), .B(n70), .Y(ab_11__16_) );
  NOR2X1 U569 ( .A(n74), .B(n70), .Y(ab_11__15_) );
  NOR2X1 U570 ( .A(n73), .B(n70), .Y(ab_11__14_) );
  NOR2X1 U571 ( .A(n72), .B(n70), .Y(ab_11__13_) );
  NOR2X1 U572 ( .A(n71), .B(n70), .Y(ab_11__12_) );
  NOR2X1 U573 ( .A(n68), .B(n70), .Y(ab_11__10_) );
  NOR2X1 U574 ( .A(n38), .B(n70), .Y(ab_11__0_) );
  NOR2X1 U575 ( .A(n67), .B(n69), .Y(ab_10__9_) );
  NOR2X1 U576 ( .A(n64), .B(n69), .Y(ab_10__8_) );
  NOR2X1 U577 ( .A(n63), .B(n69), .Y(ab_10__7_) );
  NOR2X1 U578 ( .A(n61), .B(n69), .Y(ab_10__6_) );
  NOR2X1 U579 ( .A(n60), .B(n69), .Y(ab_10__5_) );
  NOR2X1 U580 ( .A(n57), .B(n69), .Y(ab_10__4_) );
  NOR2X1 U581 ( .A(n51), .B(n69), .Y(ab_10__3_) );
  NOR2X1 U582 ( .A(n46), .B(n69), .Y(ab_10__2_) );
  NOR2X1 U583 ( .A(n81), .B(n69), .Y(ab_10__21_) );
  NOR2X1 U584 ( .A(n80), .B(n69), .Y(ab_10__20_) );
  NOR2X1 U585 ( .A(n43), .B(n69), .Y(ab_10__1_) );
  NOR2X1 U586 ( .A(n79), .B(n69), .Y(ab_10__19_) );
  NOR2X1 U587 ( .A(n78), .B(n69), .Y(ab_10__18_) );
  NOR2X1 U588 ( .A(n77), .B(n69), .Y(ab_10__17_) );
  NOR2X1 U589 ( .A(n76), .B(n69), .Y(ab_10__16_) );
  NOR2X1 U590 ( .A(n74), .B(n69), .Y(ab_10__15_) );
  NOR2X1 U591 ( .A(n73), .B(n69), .Y(ab_10__14_) );
  NOR2X1 U592 ( .A(n72), .B(n69), .Y(ab_10__13_) );
  NOR2X1 U593 ( .A(n71), .B(n69), .Y(ab_10__12_) );
  NOR2X1 U594 ( .A(n70), .B(n69), .Y(ab_10__11_) );
  NOR2X1 U595 ( .A(n38), .B(n69), .Y(ab_10__0_) );
  NOR2X1 U596 ( .A(n67), .B(n39), .Y(ab_0__9_) );
  NOR2X1 U597 ( .A(n64), .B(n39), .Y(ab_0__8_) );
  NOR2X1 U598 ( .A(n63), .B(n39), .Y(ab_0__7_) );
  NOR2X1 U599 ( .A(n61), .B(n39), .Y(ab_0__6_) );
  NOR2X1 U600 ( .A(n60), .B(n39), .Y(ab_0__5_) );
  NOR2X1 U601 ( .A(n57), .B(n39), .Y(ab_0__4_) );
  NOR2X1 U602 ( .A(n51), .B(n39), .Y(ab_0__3_) );
  NOR2X1 U603 ( .A(n75), .B(n39), .Y(ab_0__30_) );
  NOR2X1 U604 ( .A(n46), .B(n39), .Y(ab_0__2_) );
  NOR2X1 U605 ( .A(n89), .B(n38), .Y(ab_0__29_) );
  NOR2X1 U606 ( .A(n88), .B(n38), .Y(ab_0__28_) );
  NOR2X1 U607 ( .A(n87), .B(n38), .Y(ab_0__27_) );
  NOR2X1 U608 ( .A(n86), .B(n38), .Y(ab_0__26_) );
  NOR2X1 U609 ( .A(n85), .B(n38), .Y(ab_0__25_) );
  NOR2X1 U610 ( .A(n84), .B(n38), .Y(ab_0__24_) );
  NOR2X1 U611 ( .A(n83), .B(n38), .Y(ab_0__23_) );
  NOR2X1 U612 ( .A(n82), .B(n38), .Y(ab_0__22_) );
  NOR2X1 U613 ( .A(n81), .B(n38), .Y(ab_0__21_) );
  NOR2X1 U614 ( .A(n80), .B(n38), .Y(ab_0__20_) );
  NOR2X1 U615 ( .A(n43), .B(n38), .Y(ab_0__1_) );
  NOR2X1 U616 ( .A(n79), .B(n38), .Y(ab_0__19_) );
  NOR2X1 U617 ( .A(n78), .B(n38), .Y(ab_0__18_) );
  NOR2X1 U618 ( .A(n77), .B(n38), .Y(ab_0__17_) );
  NOR2X1 U619 ( .A(n76), .B(n39), .Y(ab_0__16_) );
  NOR2X1 U620 ( .A(n74), .B(n39), .Y(ab_0__15_) );
  NOR2X1 U621 ( .A(n73), .B(n39), .Y(ab_0__14_) );
  NOR2X1 U622 ( .A(n72), .B(n39), .Y(ab_0__13_) );
  NOR2X1 U623 ( .A(n71), .B(n39), .Y(ab_0__12_) );
  NOR2X1 U624 ( .A(n70), .B(n39), .Y(ab_0__11_) );
  NOR2X1 U625 ( .A(n68), .B(n39), .Y(ab_0__10_) );
endmodule


module square_root_finder_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45;
  wire   [28:13] carry;

  ADDFX2 U2_12 ( .A(A[12]), .B(n34), .CI(n1), .CO(carry[13]), .S(DIFF[12]) );
  ADDFX2 U2_13 ( .A(A[13]), .B(n33), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  ADDFX2 U2_14 ( .A(A[14]), .B(n32), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  ADDFX2 U2_15 ( .A(A[15]), .B(n31), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  ADDFX2 U2_16 ( .A(A[16]), .B(n30), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  ADDFX2 U2_17 ( .A(A[17]), .B(n29), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  ADDFX2 U2_18 ( .A(A[18]), .B(n28), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  ADDFX2 U2_19 ( .A(A[19]), .B(n27), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  ADDFX2 U2_20 ( .A(A[20]), .B(n26), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  ADDFX2 U2_21 ( .A(A[21]), .B(n25), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  ADDFX2 U2_23 ( .A(A[23]), .B(n23), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  ADDFX2 U2_27 ( .A(A[27]), .B(n19), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  ADDFX2 U2_22 ( .A(A[22]), .B(n24), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  ADDFX2 U2_24 ( .A(A[24]), .B(n22), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  ADDFX2 U2_25 ( .A(A[25]), .B(n21), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  ADDFX2 U2_26 ( .A(A[26]), .B(n20), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  AND2X2 U1 ( .A(n35), .B(n7), .Y(n1) );
  AND2X2 U2 ( .A(n42), .B(n3), .Y(n2) );
  AND2X2 U3 ( .A(n43), .B(n4), .Y(n3) );
  XOR2X1 U4 ( .A(n43), .B(n4), .Y(DIFF[3]) );
  AND2X2 U5 ( .A(n44), .B(n11), .Y(n4) );
  INVX1 U6 ( .A(B[3]), .Y(n43) );
  INVX1 U7 ( .A(B[4]), .Y(n42) );
  INVX1 U8 ( .A(B[1]), .Y(n45) );
  XOR2X1 U9 ( .A(n44), .B(n11), .Y(DIFF[2]) );
  AND2X2 U10 ( .A(n37), .B(n6), .Y(n5) );
  AND2X2 U11 ( .A(n38), .B(n9), .Y(n6) );
  AND2X2 U12 ( .A(n36), .B(n5), .Y(n7) );
  AND2X2 U13 ( .A(n40), .B(n10), .Y(n8) );
  AND2X2 U14 ( .A(n39), .B(n8), .Y(n9) );
  AND2X2 U15 ( .A(n41), .B(n2), .Y(n10) );
  AND2X2 U16 ( .A(n45), .B(n15), .Y(n11) );
  INVX1 U17 ( .A(B[2]), .Y(n44) );
  XOR2X1 U18 ( .A(n36), .B(n5), .Y(DIFF[10]) );
  XOR2X1 U19 ( .A(n37), .B(n6), .Y(DIFF[9]) );
  XOR2X1 U20 ( .A(n35), .B(n7), .Y(DIFF[11]) );
  XOR2X1 U21 ( .A(n42), .B(n3), .Y(DIFF[4]) );
  XOR2X1 U22 ( .A(n41), .B(n2), .Y(DIFF[5]) );
  XOR2X1 U23 ( .A(n40), .B(n10), .Y(DIFF[6]) );
  XOR2X1 U24 ( .A(n38), .B(n9), .Y(DIFF[8]) );
  XOR2X1 U25 ( .A(n39), .B(n8), .Y(DIFF[7]) );
  XOR2X1 U26 ( .A(n45), .B(n15), .Y(DIFF[1]) );
  INVX1 U27 ( .A(B[8]), .Y(n38) );
  INVX1 U28 ( .A(B[9]), .Y(n37) );
  INVX1 U29 ( .A(B[10]), .Y(n36) );
  INVX1 U30 ( .A(B[11]), .Y(n35) );
  INVX1 U31 ( .A(B[7]), .Y(n39) );
  INVX1 U32 ( .A(B[6]), .Y(n40) );
  INVX1 U33 ( .A(B[5]), .Y(n41) );
  INVX1 U34 ( .A(B[0]), .Y(n15) );
  XOR2X1 U35 ( .A(B[31]), .B(n14), .Y(DIFF[31]) );
  NAND2X1 U36 ( .A(n16), .B(n12), .Y(n14) );
  INVX1 U37 ( .A(B[30]), .Y(n16) );
  INVX1 U38 ( .A(B[29]), .Y(n17) );
  INVX1 U39 ( .A(B[28]), .Y(n18) );
  AND2X2 U40 ( .A(n17), .B(n13), .Y(n12) );
  XOR2X1 U41 ( .A(n18), .B(carry[28]), .Y(DIFF[28]) );
  XOR2X1 U42 ( .A(n17), .B(n13), .Y(DIFF[29]) );
  XOR2X1 U43 ( .A(n16), .B(n12), .Y(DIFF[30]) );
  AND2X2 U44 ( .A(n18), .B(carry[28]), .Y(n13) );
  INVX1 U45 ( .A(B[26]), .Y(n20) );
  INVX1 U46 ( .A(B[25]), .Y(n21) );
  INVX1 U47 ( .A(B[24]), .Y(n22) );
  INVX1 U48 ( .A(B[22]), .Y(n24) );
  INVX1 U49 ( .A(B[27]), .Y(n19) );
  INVX1 U50 ( .A(B[23]), .Y(n23) );
  INVX1 U51 ( .A(B[21]), .Y(n25) );
  INVX1 U52 ( .A(B[20]), .Y(n26) );
  INVX1 U53 ( .A(B[19]), .Y(n27) );
  INVX1 U54 ( .A(B[18]), .Y(n28) );
  INVX1 U55 ( .A(B[17]), .Y(n29) );
  INVX1 U56 ( .A(B[16]), .Y(n30) );
  INVX1 U57 ( .A(B[15]), .Y(n31) );
  INVX1 U58 ( .A(B[14]), .Y(n32) );
  INVX1 U59 ( .A(B[13]), .Y(n33) );
  INVX1 U60 ( .A(B[12]), .Y(n34) );
endmodule


module square_root_finder_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   ab_30__1_, ab_30__0_, ab_29__2_, ab_29__1_, ab_29__0_, ab_28__3_,
         ab_28__2_, ab_28__1_, ab_28__0_, ab_27__4_, ab_27__3_, ab_27__2_,
         ab_27__1_, ab_27__0_, ab_26__5_, ab_26__4_, ab_26__3_, ab_26__2_,
         ab_26__1_, ab_26__0_, ab_25__6_, ab_25__5_, ab_25__4_, ab_25__3_,
         ab_25__2_, ab_25__1_, ab_25__0_, ab_24__7_, ab_24__6_, ab_24__5_,
         ab_24__4_, ab_24__3_, ab_24__2_, ab_24__1_, ab_24__0_, ab_23__8_,
         ab_23__7_, ab_23__6_, ab_23__5_, ab_23__4_, ab_23__3_, ab_23__2_,
         ab_23__1_, ab_23__0_, ab_22__9_, ab_22__8_, ab_22__7_, ab_22__6_,
         ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_, ab_22__0_,
         ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_, ab_21__6_, ab_21__5_,
         ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_, ab_21__0_, ab_20__11_,
         ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_, ab_20__6_, ab_20__5_,
         ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_, ab_20__0_, ab_19__12_,
         ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_, ab_19__6_,
         ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_, ab_19__0_,
         ab_18__13_, ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_, ab_18__8_,
         ab_18__7_, ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_, ab_18__2_,
         ab_18__1_, ab_18__0_, ab_17__14_, ab_17__13_, ab_17__12_, ab_17__11_,
         ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_, ab_17__6_, ab_17__5_,
         ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_, ab_17__0_, ab_16__15_,
         ab_16__14_, ab_16__13_, ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_,
         ab_16__8_, ab_16__7_, ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_,
         ab_16__2_, ab_16__1_, ab_16__0_, ab_15__16_, ab_15__14_, ab_15__13_,
         ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_,
         ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_,
         ab_15__0_, ab_14__17_, ab_14__16_, ab_14__15_, ab_14__13_, ab_14__12_,
         ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_, ab_14__6_,
         ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_, ab_14__0_,
         ab_13__18_, ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_,
         ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_,
         ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_,
         ab_13__0_, ab_12__19_, ab_12__18_, ab_12__17_, ab_12__16_, ab_12__15_,
         ab_12__14_, ab_12__13_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_,
         ab_12__7_, ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_,
         ab_12__1_, ab_12__0_, ab_11__20_, ab_11__19_, ab_11__18_, ab_11__17_,
         ab_11__16_, ab_11__15_, ab_11__14_, ab_11__13_, ab_11__12_,
         ab_11__10_, ab_11__9_, ab_11__8_, ab_11__7_, ab_11__6_, ab_11__5_,
         ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_, ab_11__0_, ab_10__21_,
         ab_10__20_, ab_10__19_, ab_10__18_, ab_10__17_, ab_10__16_,
         ab_10__15_, ab_10__14_, ab_10__13_, ab_10__12_, ab_10__11_, ab_10__9_,
         ab_10__8_, ab_10__7_, ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_,
         ab_10__2_, ab_10__1_, ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_,
         ab_9__19_, ab_9__18_, ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_,
         ab_9__13_, ab_9__12_, ab_9__11_, ab_9__10_, ab_9__8_, ab_9__7_,
         ab_9__6_, ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_,
         ab_8__23_, ab_8__22_, ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_,
         ab_8__17_, ab_8__16_, ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_,
         ab_8__11_, ab_8__10_, ab_8__9_, ab_8__7_, ab_8__6_, ab_8__5_,
         ab_8__4_, ab_8__3_, ab_8__2_, ab_8__1_, ab_8__0_, ab_7__24_,
         ab_7__23_, ab_7__22_, ab_7__21_, ab_7__20_, ab_7__19_, ab_7__18_,
         ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_, ab_7__13_, ab_7__12_,
         ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_, ab_7__6_, ab_7__5_,
         ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_, ab_7__0_, ab_6__25_,
         ab_6__24_, ab_6__23_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_,
         ab_6__18_, ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_,
         ab_6__12_, ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__26_,
         ab_5__25_, ab_5__24_, ab_5__23_, ab_5__22_, ab_5__21_, ab_5__20_,
         ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_, ab_5__15_, ab_5__14_,
         ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_, ab_5__9_, ab_5__8_,
         ab_5__7_, ab_5__6_, ab_5__4_, ab_5__3_, ab_5__2_, ab_5__1_, ab_5__0_,
         ab_4__27_, ab_4__26_, ab_4__25_, ab_4__24_, ab_4__23_, ab_4__22_,
         ab_4__21_, ab_4__20_, ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_,
         ab_4__15_, ab_4__14_, ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_,
         ab_4__9_, ab_4__8_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__3_, ab_4__2_,
         ab_4__1_, ab_4__0_, ab_3__28_, ab_3__27_, ab_3__26_, ab_3__25_,
         ab_3__24_, ab_3__23_, ab_3__22_, ab_3__21_, ab_3__20_, ab_3__19_,
         ab_3__18_, ab_3__17_, ab_3__16_, ab_3__15_, ab_3__14_, ab_3__13_,
         ab_3__12_, ab_3__11_, ab_3__10_, ab_3__9_, ab_3__8_, ab_3__7_,
         ab_3__6_, ab_3__5_, ab_3__4_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__29_,
         ab_2__28_, ab_2__27_, ab_2__26_, ab_2__25_, ab_2__24_, ab_2__23_,
         ab_2__22_, ab_2__21_, ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_,
         ab_2__16_, ab_2__15_, ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_,
         ab_2__10_, ab_2__9_, ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_,
         ab_2__3_, ab_2__1_, ab_2__0_, ab_1__30_, ab_1__29_, ab_1__28_,
         ab_1__27_, ab_1__26_, ab_1__25_, ab_1__24_, ab_1__23_, ab_1__22_,
         ab_1__21_, ab_1__20_, ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_,
         ab_1__15_, ab_1__14_, ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_,
         ab_1__9_, ab_1__8_, ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_,
         ab_1__2_, ab_1__0_, ab_0__30_, ab_0__29_, ab_0__28_, ab_0__27_,
         ab_0__26_, ab_0__25_, ab_0__24_, ab_0__23_, ab_0__22_, ab_0__21_,
         ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_, ab_0__16_, ab_0__15_,
         ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_, ab_0__10_, ab_0__9_,
         ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_,
         ab_0__1_, CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_,
         CARRYB_15__12_, CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_,
         CARRYB_15__8_, CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_,
         CARRYB_15__4_, CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_,
         CARRYB_15__0_, CARRYB_14__16_, CARRYB_14__15_, CARRYB_14__14_,
         CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_, CARRYB_14__10_,
         CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_, CARRYB_14__6_,
         CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_, CARRYB_14__2_,
         CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__17_, CARRYB_13__16_,
         CARRYB_13__15_, CARRYB_13__14_, CARRYB_13__13_, CARRYB_13__12_,
         CARRYB_13__11_, CARRYB_13__10_, CARRYB_13__9_, CARRYB_13__8_,
         CARRYB_13__7_, CARRYB_13__6_, CARRYB_13__5_, CARRYB_13__4_,
         CARRYB_13__3_, CARRYB_13__2_, CARRYB_13__1_, CARRYB_13__0_,
         CARRYB_12__18_, CARRYB_12__17_, CARRYB_12__16_, CARRYB_12__15_,
         CARRYB_12__14_, CARRYB_12__13_, CARRYB_12__12_, CARRYB_12__11_,
         CARRYB_12__10_, CARRYB_12__9_, CARRYB_12__8_, CARRYB_12__7_,
         CARRYB_12__6_, CARRYB_12__5_, CARRYB_12__4_, CARRYB_12__3_,
         CARRYB_12__2_, CARRYB_12__1_, CARRYB_12__0_, CARRYB_11__19_,
         CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_, CARRYB_11__15_,
         CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_, CARRYB_11__11_,
         CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_, CARRYB_11__7_,
         CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_, CARRYB_11__3_,
         CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_, CARRYB_10__20_,
         CARRYB_10__19_, CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_,
         CARRYB_10__15_, CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_,
         CARRYB_10__11_, CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_,
         CARRYB_10__7_, CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_,
         CARRYB_10__3_, CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__23_, CARRYB_7__22_, CARRYB_7__21_,
         CARRYB_7__20_, CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_,
         CARRYB_7__16_, CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_,
         CARRYB_7__12_, CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_,
         CARRYB_7__8_, CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_,
         CARRYB_7__3_, CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__24_,
         CARRYB_6__23_, CARRYB_6__22_, CARRYB_6__21_, CARRYB_6__20_,
         CARRYB_6__19_, CARRYB_6__18_, CARRYB_6__17_, CARRYB_6__16_,
         CARRYB_6__15_, CARRYB_6__14_, CARRYB_6__13_, CARRYB_6__12_,
         CARRYB_6__11_, CARRYB_6__10_, CARRYB_6__9_, CARRYB_6__8_,
         CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_, CARRYB_6__4_, CARRYB_6__3_,
         CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_, CARRYB_5__25_,
         CARRYB_5__24_, CARRYB_5__23_, CARRYB_5__22_, CARRYB_5__21_,
         CARRYB_5__20_, CARRYB_5__19_, CARRYB_5__18_, CARRYB_5__17_,
         CARRYB_5__16_, CARRYB_5__15_, CARRYB_5__14_, CARRYB_5__13_,
         CARRYB_5__12_, CARRYB_5__11_, CARRYB_5__10_, CARRYB_5__9_,
         CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_,
         CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__26_,
         CARRYB_4__25_, CARRYB_4__24_, CARRYB_4__23_, CARRYB_4__22_,
         CARRYB_4__21_, CARRYB_4__20_, CARRYB_4__19_, CARRYB_4__18_,
         CARRYB_4__17_, CARRYB_4__16_, CARRYB_4__15_, CARRYB_4__14_,
         CARRYB_4__13_, CARRYB_4__12_, CARRYB_4__11_, CARRYB_4__10_,
         CARRYB_4__9_, CARRYB_4__8_, CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_,
         CARRYB_4__4_, CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_,
         CARRYB_3__27_, CARRYB_3__26_, CARRYB_3__25_, CARRYB_3__24_,
         CARRYB_3__23_, CARRYB_3__22_, CARRYB_3__21_, CARRYB_3__20_,
         CARRYB_3__19_, CARRYB_3__18_, CARRYB_3__17_, CARRYB_3__16_,
         CARRYB_3__15_, CARRYB_3__14_, CARRYB_3__13_, CARRYB_3__12_,
         CARRYB_3__11_, CARRYB_3__10_, CARRYB_3__9_, CARRYB_3__8_,
         CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_,
         CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_, CARRYB_2__28_,
         CARRYB_2__27_, CARRYB_2__26_, CARRYB_2__25_, CARRYB_2__24_,
         CARRYB_2__23_, CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_,
         CARRYB_2__19_, CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_,
         CARRYB_2__15_, CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_,
         CARRYB_2__11_, CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_,
         CARRYB_2__7_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_15__16_, SUMB_15__15_,
         SUMB_15__14_, SUMB_15__13_, SUMB_15__12_, SUMB_15__11_, SUMB_15__10_,
         SUMB_15__9_, SUMB_15__8_, SUMB_15__7_, SUMB_15__6_, SUMB_15__5_,
         SUMB_15__4_, SUMB_15__3_, SUMB_15__2_, SUMB_15__1_, SUMB_14__17_,
         SUMB_14__16_, SUMB_14__15_, SUMB_14__14_, SUMB_14__13_, SUMB_14__12_,
         SUMB_14__11_, SUMB_14__10_, SUMB_14__9_, SUMB_14__8_, SUMB_14__7_,
         SUMB_14__6_, SUMB_14__5_, SUMB_14__4_, SUMB_14__3_, SUMB_14__2_,
         SUMB_14__1_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_, SUMB_13__15_,
         SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_, SUMB_13__10_,
         SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_, SUMB_13__5_,
         SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_, SUMB_12__19_,
         SUMB_12__18_, SUMB_12__17_, SUMB_12__16_, SUMB_12__15_, SUMB_12__14_,
         SUMB_12__13_, SUMB_12__12_, SUMB_12__11_, SUMB_12__10_, SUMB_12__9_,
         SUMB_12__8_, SUMB_12__7_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_,
         SUMB_12__3_, SUMB_12__2_, SUMB_12__1_, SUMB_11__20_, SUMB_11__19_,
         SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_, SUMB_11__14_,
         SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_, SUMB_11__9_,
         SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_, SUMB_11__4_,
         SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__21_, SUMB_10__20_,
         SUMB_10__19_, SUMB_10__18_, SUMB_10__17_, SUMB_10__16_, SUMB_10__15_,
         SUMB_10__14_, SUMB_10__13_, SUMB_10__12_, SUMB_10__11_, SUMB_10__10_,
         SUMB_10__9_, SUMB_10__8_, SUMB_10__7_, SUMB_10__6_, SUMB_10__5_,
         SUMB_10__4_, SUMB_10__3_, SUMB_10__2_, SUMB_10__1_, SUMB_9__22_,
         SUMB_9__21_, SUMB_9__20_, SUMB_9__19_, SUMB_9__18_, SUMB_9__17_,
         SUMB_9__16_, SUMB_9__15_, SUMB_9__14_, SUMB_9__13_, SUMB_9__12_,
         SUMB_9__11_, SUMB_9__10_, SUMB_9__9_, SUMB_9__8_, SUMB_9__7_,
         SUMB_9__6_, SUMB_9__5_, SUMB_9__4_, SUMB_9__3_, SUMB_9__2_,
         SUMB_9__1_, SUMB_8__23_, SUMB_8__22_, SUMB_8__21_, SUMB_8__20_,
         SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_, SUMB_8__15_,
         SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_, SUMB_8__10_,
         SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_, SUMB_8__5_,
         SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_, SUMB_7__24_,
         SUMB_7__23_, SUMB_7__22_, SUMB_7__21_, SUMB_7__20_, SUMB_7__19_,
         SUMB_7__18_, SUMB_7__17_, SUMB_7__16_, SUMB_7__15_, SUMB_7__14_,
         SUMB_7__13_, SUMB_7__12_, SUMB_7__11_, SUMB_7__10_, SUMB_7__9_,
         SUMB_7__8_, SUMB_7__7_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_,
         SUMB_7__3_, SUMB_7__2_, SUMB_7__1_, SUMB_6__25_, SUMB_6__24_,
         SUMB_6__23_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_, SUMB_6__19_,
         SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_, SUMB_6__14_,
         SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_, SUMB_6__9_,
         SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_,
         SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__26_, SUMB_5__25_,
         SUMB_5__24_, SUMB_5__23_, SUMB_5__22_, SUMB_5__21_, SUMB_5__20_,
         SUMB_5__19_, SUMB_5__18_, SUMB_5__17_, SUMB_5__16_, SUMB_5__15_,
         SUMB_5__14_, SUMB_5__13_, SUMB_5__12_, SUMB_5__11_, SUMB_5__10_,
         SUMB_5__9_, SUMB_5__8_, SUMB_5__7_, SUMB_5__6_, SUMB_5__5_,
         SUMB_5__4_, SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__27_,
         SUMB_4__26_, SUMB_4__25_, SUMB_4__24_, SUMB_4__23_, SUMB_4__22_,
         SUMB_4__21_, SUMB_4__20_, SUMB_4__19_, SUMB_4__18_, SUMB_4__17_,
         SUMB_4__16_, SUMB_4__15_, SUMB_4__14_, SUMB_4__13_, SUMB_4__12_,
         SUMB_4__11_, SUMB_4__10_, SUMB_4__9_, SUMB_4__8_, SUMB_4__7_,
         SUMB_4__6_, SUMB_4__5_, SUMB_4__4_, SUMB_4__3_, SUMB_4__2_,
         SUMB_4__1_, SUMB_3__28_, SUMB_3__27_, SUMB_3__26_, SUMB_3__25_,
         SUMB_3__24_, SUMB_3__23_, SUMB_3__22_, SUMB_3__21_, SUMB_3__20_,
         SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_, SUMB_3__15_,
         SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_, SUMB_3__10_,
         SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_, SUMB_3__5_,
         SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_, SUMB_2__29_,
         SUMB_2__28_, SUMB_2__27_, SUMB_2__26_, SUMB_2__25_, SUMB_2__24_,
         SUMB_2__23_, SUMB_2__22_, SUMB_2__21_, SUMB_2__20_, SUMB_2__19_,
         SUMB_2__18_, SUMB_2__17_, SUMB_2__16_, SUMB_2__15_, SUMB_2__14_,
         SUMB_2__13_, SUMB_2__12_, SUMB_2__11_, SUMB_2__10_, SUMB_2__9_,
         SUMB_2__8_, SUMB_2__7_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_,
         SUMB_2__3_, SUMB_2__2_, SUMB_2__1_, SUMB_1__29_, SUMB_1__28_,
         SUMB_1__27_, SUMB_1__26_, SUMB_1__25_, SUMB_1__24_, SUMB_1__23_,
         SUMB_1__22_, SUMB_1__21_, SUMB_1__20_, SUMB_1__19_, SUMB_1__18_,
         SUMB_1__17_, SUMB_1__16_, SUMB_1__15_, SUMB_1__14_, SUMB_1__13_,
         SUMB_1__12_, SUMB_1__11_, SUMB_1__10_, SUMB_1__9_, SUMB_1__8_,
         SUMB_1__7_, SUMB_1__6_, SUMB_1__5_, SUMB_1__4_, SUMB_1__3_,
         SUMB_1__2_, SUMB_1__1_, CARRYB_30__0_, CARRYB_29__1_, CARRYB_29__0_,
         CARRYB_28__2_, CARRYB_28__1_, CARRYB_28__0_, CARRYB_27__3_,
         CARRYB_27__2_, CARRYB_27__1_, CARRYB_27__0_, CARRYB_26__4_,
         CARRYB_26__3_, CARRYB_26__2_, CARRYB_26__1_, CARRYB_26__0_,
         CARRYB_25__5_, CARRYB_25__4_, CARRYB_25__3_, CARRYB_25__2_,
         CARRYB_25__1_, CARRYB_25__0_, CARRYB_24__6_, CARRYB_24__5_,
         CARRYB_24__4_, CARRYB_24__3_, CARRYB_24__2_, CARRYB_24__1_,
         CARRYB_24__0_, CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_,
         CARRYB_23__4_, CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_,
         CARRYB_23__0_, CARRYB_22__8_, CARRYB_22__7_, CARRYB_22__6_,
         CARRYB_22__5_, CARRYB_22__4_, CARRYB_22__3_, CARRYB_22__2_,
         CARRYB_22__1_, CARRYB_22__0_, CARRYB_21__9_, CARRYB_21__8_,
         CARRYB_21__7_, CARRYB_21__6_, CARRYB_21__5_, CARRYB_21__4_,
         CARRYB_21__3_, CARRYB_21__2_, CARRYB_21__1_, CARRYB_21__0_,
         CARRYB_20__10_, CARRYB_20__9_, CARRYB_20__8_, CARRYB_20__7_,
         CARRYB_20__6_, CARRYB_20__5_, CARRYB_20__4_, CARRYB_20__3_,
         CARRYB_20__2_, CARRYB_20__1_, CARRYB_20__0_, CARRYB_19__11_,
         CARRYB_19__10_, CARRYB_19__9_, CARRYB_19__8_, CARRYB_19__7_,
         CARRYB_19__6_, CARRYB_19__5_, CARRYB_19__4_, CARRYB_19__3_,
         CARRYB_19__2_, CARRYB_19__1_, CARRYB_19__0_, CARRYB_18__12_,
         CARRYB_18__11_, CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_,
         CARRYB_18__7_, CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_,
         CARRYB_18__3_, CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_,
         CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_, CARRYB_17__10_,
         CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_, CARRYB_17__6_,
         CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_, CARRYB_17__2_,
         CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__14_, CARRYB_16__13_,
         CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_, CARRYB_16__9_,
         CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_, CARRYB_16__5_,
         CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_,
         CARRYB_16__0_, SUMB_30__1_, SUMB_29__2_, SUMB_29__1_, SUMB_28__3_,
         SUMB_28__2_, SUMB_28__1_, SUMB_27__4_, SUMB_27__3_, SUMB_27__2_,
         SUMB_27__1_, SUMB_26__5_, SUMB_26__4_, SUMB_26__3_, SUMB_26__2_,
         SUMB_26__1_, SUMB_25__6_, SUMB_25__5_, SUMB_25__4_, SUMB_25__3_,
         SUMB_25__2_, SUMB_25__1_, SUMB_24__7_, SUMB_24__6_, SUMB_24__5_,
         SUMB_24__4_, SUMB_24__3_, SUMB_24__2_, SUMB_24__1_, SUMB_23__8_,
         SUMB_23__7_, SUMB_23__6_, SUMB_23__5_, SUMB_23__4_, SUMB_23__3_,
         SUMB_23__2_, SUMB_23__1_, SUMB_22__9_, SUMB_22__8_, SUMB_22__7_,
         SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_, SUMB_22__2_,
         SUMB_22__1_, SUMB_21__10_, SUMB_21__9_, SUMB_21__8_, SUMB_21__7_,
         SUMB_21__6_, SUMB_21__5_, SUMB_21__4_, SUMB_21__3_, SUMB_21__2_,
         SUMB_21__1_, SUMB_20__11_, SUMB_20__10_, SUMB_20__9_, SUMB_20__8_,
         SUMB_20__7_, SUMB_20__6_, SUMB_20__5_, SUMB_20__4_, SUMB_20__3_,
         SUMB_20__2_, SUMB_20__1_, SUMB_19__12_, SUMB_19__11_, SUMB_19__10_,
         SUMB_19__9_, SUMB_19__8_, SUMB_19__7_, SUMB_19__6_, SUMB_19__5_,
         SUMB_19__4_, SUMB_19__3_, SUMB_19__2_, SUMB_19__1_, SUMB_18__13_,
         SUMB_18__12_, SUMB_18__11_, SUMB_18__10_, SUMB_18__9_, SUMB_18__8_,
         SUMB_18__7_, SUMB_18__6_, SUMB_18__5_, SUMB_18__4_, SUMB_18__3_,
         SUMB_18__2_, SUMB_18__1_, SUMB_17__14_, SUMB_17__13_, SUMB_17__12_,
         SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_, SUMB_17__7_,
         SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_, SUMB_17__2_,
         SUMB_17__1_, SUMB_16__15_, SUMB_16__14_, SUMB_16__13_, SUMB_16__12_,
         SUMB_16__11_, SUMB_16__10_, SUMB_16__9_, SUMB_16__8_, SUMB_16__7_,
         SUMB_16__6_, SUMB_16__5_, SUMB_16__4_, SUMB_16__3_, SUMB_16__2_,
         SUMB_16__1_, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82;

  ADDFX2 S2_2_28 ( .A(ab_2__28_), .B(n35), .CI(SUMB_1__29_), .CO(CARRYB_2__28_), .S(SUMB_2__28_) );
  ADDFX2 S2_2_27 ( .A(ab_2__27_), .B(n34), .CI(SUMB_1__28_), .CO(CARRYB_2__27_), .S(SUMB_2__27_) );
  ADDFX2 S2_2_26 ( .A(ab_2__26_), .B(n33), .CI(SUMB_1__27_), .CO(CARRYB_2__26_), .S(SUMB_2__26_) );
  ADDFX2 S2_2_25 ( .A(ab_2__25_), .B(n32), .CI(SUMB_1__26_), .CO(CARRYB_2__25_), .S(SUMB_2__25_) );
  ADDFX2 S2_2_24 ( .A(ab_2__24_), .B(n31), .CI(SUMB_1__25_), .CO(CARRYB_2__24_), .S(SUMB_2__24_) );
  ADDFX2 S2_2_23 ( .A(ab_2__23_), .B(n30), .CI(SUMB_1__24_), .CO(CARRYB_2__23_), .S(SUMB_2__23_) );
  ADDFX2 S2_2_22 ( .A(ab_2__22_), .B(n29), .CI(SUMB_1__23_), .CO(CARRYB_2__22_), .S(SUMB_2__22_) );
  ADDFX2 S2_2_21 ( .A(ab_2__21_), .B(n28), .CI(SUMB_1__22_), .CO(CARRYB_2__21_), .S(SUMB_2__21_) );
  ADDFX2 S2_2_20 ( .A(ab_2__20_), .B(n27), .CI(SUMB_1__21_), .CO(CARRYB_2__20_), .S(SUMB_2__20_) );
  ADDFX2 S2_2_19 ( .A(ab_2__19_), .B(n26), .CI(SUMB_1__20_), .CO(CARRYB_2__19_), .S(SUMB_2__19_) );
  ADDFX2 S2_2_18 ( .A(ab_2__18_), .B(n25), .CI(SUMB_1__19_), .CO(CARRYB_2__18_), .S(SUMB_2__18_) );
  ADDFX2 S2_2_17 ( .A(ab_2__17_), .B(n24), .CI(SUMB_1__18_), .CO(CARRYB_2__17_), .S(SUMB_2__17_) );
  ADDFX2 S2_2_16 ( .A(ab_2__16_), .B(n23), .CI(SUMB_1__17_), .CO(CARRYB_2__16_), .S(SUMB_2__16_) );
  XOR3X2 S2_23_8 ( .A(ab_23__8_), .B(CARRYB_22__8_), .C(SUMB_22__9_), .Y(
        SUMB_23__8_) );
  XOR3X2 S2_24_7 ( .A(ab_24__7_), .B(CARRYB_23__7_), .C(SUMB_23__8_), .Y(
        SUMB_24__7_) );
  XOR3X2 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .C(SUMB_20__11_), .Y(
        SUMB_21__10_) );
  XOR3X2 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .C(SUMB_21__10_), .Y(
        SUMB_22__9_) );
  XOR3X2 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .C(SUMB_18__13_), .Y(
        SUMB_19__12_) );
  XOR3X2 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .C(SUMB_19__12_), .Y(
        SUMB_20__11_) );
  XOR3X2 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .C(SUMB_16__15_), .Y(
        SUMB_17__14_) );
  XOR3X2 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .C(SUMB_17__14_), .Y(
        SUMB_18__13_) );
  XOR3X2 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .C(SUMB_14__17_), .Y(
        SUMB_15__16_) );
  XOR3X2 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .C(SUMB_15__16_), .Y(
        SUMB_16__15_) );
  XOR3X2 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .C(SUMB_12__19_), .Y(
        SUMB_13__18_) );
  XOR3X2 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .C(SUMB_13__18_), .Y(
        SUMB_14__17_) );
  XOR3X2 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .C(SUMB_10__21_), .Y(
        SUMB_11__20_) );
  XOR3X2 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .C(SUMB_11__20_), .Y(
        SUMB_12__19_) );
  XOR3X2 S2_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .C(SUMB_8__23_), .Y(
        SUMB_9__22_) );
  XOR3X2 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .C(SUMB_9__22_), .Y(
        SUMB_10__21_) );
  XOR3X2 S2_7_24 ( .A(ab_7__24_), .B(CARRYB_6__24_), .C(SUMB_6__25_), .Y(
        SUMB_7__24_) );
  XOR3X2 S2_8_23 ( .A(ab_8__23_), .B(CARRYB_7__23_), .C(SUMB_7__24_), .Y(
        SUMB_8__23_) );
  XOR3X2 S2_5_26 ( .A(ab_5__26_), .B(CARRYB_4__26_), .C(SUMB_4__27_), .Y(
        SUMB_5__26_) );
  XOR3X2 S2_6_25 ( .A(ab_6__25_), .B(CARRYB_5__25_), .C(SUMB_5__26_), .Y(
        SUMB_6__25_) );
  XOR3X2 S2_3_28 ( .A(ab_3__28_), .B(CARRYB_2__28_), .C(SUMB_2__29_), .Y(
        SUMB_3__28_) );
  XOR3X2 S2_4_27 ( .A(ab_4__27_), .B(CARRYB_3__27_), .C(SUMB_3__28_), .Y(
        SUMB_4__27_) );
  ADDFX2 S2_3_27 ( .A(ab_3__27_), .B(CARRYB_2__27_), .CI(SUMB_2__28_), .CO(
        CARRYB_3__27_), .S(SUMB_3__27_) );
  ADDFX2 S2_3_24 ( .A(ab_3__24_), .B(CARRYB_2__24_), .CI(SUMB_2__25_), .CO(
        CARRYB_3__24_), .S(SUMB_3__24_) );
  XOR3X2 S2_2_29 ( .A(ab_2__29_), .B(n36), .C(ab_1__30_), .Y(SUMB_2__29_) );
  ADDFX2 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  ADDFX2 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  ADDFX2 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), 
        .CO(CARRYB_20__10_), .S(SUMB_20__10_) );
  ADDFX2 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  ADDFX2 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  ADDFX2 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), 
        .CO(CARRYB_18__12_), .S(SUMB_18__12_) );
  ADDFX2 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), 
        .CO(CARRYB_18__11_), .S(SUMB_18__11_) );
  ADDFX2 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), 
        .CO(CARRYB_18__10_), .S(SUMB_18__10_) );
  ADDFX2 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  ADDFX2 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  ADDFX2 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  ADDFX2 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), 
        .CO(CARRYB_12__18_), .S(SUMB_12__18_) );
  ADDFX2 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), 
        .CO(CARRYB_12__17_), .S(SUMB_12__17_) );
  ADDFX2 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), 
        .CO(CARRYB_12__16_), .S(SUMB_12__16_) );
  ADDFX2 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), 
        .CO(CARRYB_11__16_), .S(SUMB_11__16_) );
  ADDFX2 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  ADDFX2 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  ADDFX2 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  ADDFX2 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  ADDFX2 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  ADDFX2 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  ADDFX2 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  ADDFX2 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  ADDFX2 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), 
        .CO(CARRYB_19__11_), .S(SUMB_19__11_) );
  ADDFX2 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), 
        .CO(CARRYB_19__10_), .S(SUMB_19__10_) );
  ADDFX2 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  ADDFX2 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  ADDFX2 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  ADDFX2 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), 
        .CO(CARRYB_17__13_), .S(SUMB_17__13_) );
  ADDFX2 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), 
        .CO(CARRYB_17__12_), .S(SUMB_17__12_) );
  ADDFX2 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  ADDFX2 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  ADDFX2 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  ADDFX2 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  ADDFX2 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), 
        .CO(CARRYB_14__16_), .S(SUMB_14__16_) );
  ADDFX2 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), 
        .CO(CARRYB_13__17_), .S(SUMB_13__17_) );
  ADDFX2 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), 
        .CO(CARRYB_13__16_), .S(SUMB_13__16_) );
  ADDFX2 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), 
        .CO(CARRYB_11__19_), .S(SUMB_11__19_) );
  ADDFX2 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), 
        .CO(CARRYB_11__17_), .S(SUMB_11__17_) );
  ADDFX2 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  ADDFX2 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), 
        .CO(CARRYB_17__11_), .S(SUMB_17__11_) );
  ADDFX2 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), 
        .CO(CARRYB_17__10_), .S(SUMB_17__10_) );
  ADDFX2 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  ADDFX2 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  ADDFX2 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), 
        .CO(CARRYB_16__14_), .S(SUMB_16__14_) );
  ADDFX2 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), 
        .CO(CARRYB_16__13_), .S(SUMB_16__13_) );
  ADDFX2 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), 
        .CO(CARRYB_16__12_), .S(SUMB_16__12_) );
  ADDFX2 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), 
        .CO(CARRYB_16__11_), .S(SUMB_16__11_) );
  ADDFX2 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), 
        .CO(CARRYB_16__10_), .S(SUMB_16__10_) );
  ADDFX2 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), 
        .CO(CARRYB_11__18_), .S(SUMB_11__18_) );
  ADDFX2 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  ADDFX2 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  ADDFX2 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  ADDFX2 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  ADDFX2 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  ADDFX2 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  ADDFX2 S2_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(SUMB_7__23_), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  ADDFX2 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  ADDFX2 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  ADDFX2 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  ADDFX2 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  ADDFX2 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  ADDFX2 S2_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(SUMB_6__23_), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  ADDFX2 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  ADDFX2 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  ADDFX2 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  ADDFX2 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  ADDFX2 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  ADDFX2 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  ADDFX2 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  ADDFX2 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  ADDFX2 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  ADDFX2 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  ADDFX2 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  ADDFX2 S2_5_24 ( .A(ab_5__24_), .B(CARRYB_4__24_), .CI(SUMB_4__25_), .CO(
        CARRYB_5__24_), .S(SUMB_5__24_) );
  ADDFX2 S2_5_23 ( .A(ab_5__23_), .B(CARRYB_4__23_), .CI(SUMB_4__24_), .CO(
        CARRYB_5__23_), .S(SUMB_5__23_) );
  ADDFX2 S2_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(SUMB_4__23_), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  ADDFX2 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  ADDFX2 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  ADDFX2 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  ADDFX2 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  ADDFX2 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  ADDFX2 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  ADDFX2 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  ADDFX2 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  ADDFX2 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  ADDFX2 S2_3_25 ( .A(ab_3__25_), .B(CARRYB_2__25_), .CI(SUMB_2__26_), .CO(
        CARRYB_3__25_), .S(SUMB_3__25_) );
  ADDFX2 S2_3_23 ( .A(ab_3__23_), .B(CARRYB_2__23_), .CI(SUMB_2__24_), .CO(
        CARRYB_3__23_), .S(SUMB_3__23_) );
  ADDFX2 S2_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(SUMB_2__23_), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  ADDFX2 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  ADDFX2 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  ADDFX2 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  ADDFX2 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  ADDFX2 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  ADDFX2 S2_23_7 ( .A(ab_23__7_), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  ADDFX2 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  ADDFX2 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  ADDFX2 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  ADDFX2 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  ADDFX2 S2_7_23 ( .A(ab_7__23_), .B(CARRYB_6__23_), .CI(SUMB_6__24_), .CO(
        CARRYB_7__23_), .S(SUMB_7__23_) );
  ADDFX2 S2_6_24 ( .A(ab_6__24_), .B(CARRYB_5__24_), .CI(SUMB_5__25_), .CO(
        CARRYB_6__24_), .S(SUMB_6__24_) );
  ADDFX2 S2_6_23 ( .A(ab_6__23_), .B(CARRYB_5__23_), .CI(SUMB_5__24_), .CO(
        CARRYB_6__23_), .S(SUMB_6__23_) );
  ADDFX2 S2_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(SUMB_5__23_), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  ADDFX2 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  ADDFX2 S2_5_25 ( .A(ab_5__25_), .B(CARRYB_4__25_), .CI(SUMB_4__26_), .CO(
        CARRYB_5__25_), .S(SUMB_5__25_) );
  ADDFX2 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  ADDFX2 S2_4_26 ( .A(ab_4__26_), .B(CARRYB_3__26_), .CI(SUMB_3__27_), .CO(
        CARRYB_4__26_), .S(SUMB_4__26_) );
  ADDFX2 S2_4_25 ( .A(ab_4__25_), .B(CARRYB_3__25_), .CI(SUMB_3__26_), .CO(
        CARRYB_4__25_), .S(SUMB_4__25_) );
  ADDFX2 S2_4_24 ( .A(ab_4__24_), .B(CARRYB_3__24_), .CI(SUMB_3__25_), .CO(
        CARRYB_4__24_), .S(SUMB_4__24_) );
  ADDFX2 S2_4_23 ( .A(ab_4__23_), .B(CARRYB_3__23_), .CI(SUMB_3__24_), .CO(
        CARRYB_4__23_), .S(SUMB_4__23_) );
  ADDFX2 S2_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(SUMB_3__23_), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  ADDFX2 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  ADDFX2 S2_3_26 ( .A(ab_3__26_), .B(CARRYB_2__26_), .CI(SUMB_2__27_), .CO(
        CARRYB_3__26_), .S(SUMB_3__26_) );
  ADDFX2 S2_12_12 ( .A(B[12]), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  ADDFX2 S2_15_15 ( .A(B[15]), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  ADDFX2 S2_14_14 ( .A(B[14]), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  ADDFX2 S2_13_13 ( .A(B[13]), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  ADDFX2 S2_11_11 ( .A(B[11]), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  ADDFX2 S2_10_10 ( .A(B[10]), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  ADDFX2 S2_9_9 ( .A(B[9]), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  ADDFX2 S2_8_8 ( .A(B[8]), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  ADDFX2 S2_7_7 ( .A(B[7]), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  XOR3X2 S2_27_4 ( .A(ab_27__4_), .B(CARRYB_26__4_), .C(SUMB_26__5_), .Y(
        SUMB_27__4_) );
  XOR3X2 S2_28_3 ( .A(ab_28__3_), .B(CARRYB_27__3_), .C(SUMB_27__4_), .Y(
        SUMB_28__3_) );
  XOR3X2 S2_25_6 ( .A(ab_25__6_), .B(CARRYB_24__6_), .C(SUMB_24__7_), .Y(
        SUMB_25__6_) );
  XOR3X2 S2_26_5 ( .A(ab_26__5_), .B(CARRYB_25__5_), .C(SUMB_25__6_), .Y(
        SUMB_26__5_) );
  ADDFX2 S1_30_0 ( .A(ab_30__0_), .B(CARRYB_29__0_), .CI(SUMB_29__1_), .CO(
        CARRYB_30__0_), .S(PRODUCT[30]) );
  ADDFX2 S1_29_0 ( .A(ab_29__0_), .B(CARRYB_28__0_), .CI(SUMB_28__1_), .CO(
        CARRYB_29__0_), .S(PRODUCT[29]) );
  ADDFX2 S1_28_0 ( .A(ab_28__0_), .B(CARRYB_27__0_), .CI(SUMB_27__1_), .CO(
        CARRYB_28__0_), .S(PRODUCT[28]) );
  ADDFX2 S2_29_1 ( .A(ab_29__1_), .B(CARRYB_28__1_), .CI(SUMB_28__2_), .CO(
        CARRYB_29__1_), .S(SUMB_29__1_) );
  ADDFX2 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(PRODUCT[18]) );
  ADDFX2 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  ADDFX2 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  ADDFX2 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  ADDFX2 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  ADDFX2 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  ADDFX2 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  ADDFX2 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(PRODUCT[17]) );
  ADDFX2 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(PRODUCT[16]) );
  ADDFX2 S1_26_0 ( .A(ab_26__0_), .B(CARRYB_25__0_), .CI(SUMB_25__1_), .CO(
        CARRYB_26__0_), .S(PRODUCT[26]) );
  ADDFX2 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  ADDFX2 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  ADDFX2 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  ADDFX2 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  ADDFX2 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  ADDFX2 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  ADDFX2 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  ADDFX2 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  ADDFX2 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  ADDFX2 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  ADDFX2 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  ADDFX2 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  ADDFX2 S1_27_0 ( .A(ab_27__0_), .B(CARRYB_26__0_), .CI(SUMB_26__1_), .CO(
        CARRYB_27__0_), .S(PRODUCT[27]) );
  ADDFX2 S2_28_2 ( .A(ab_28__2_), .B(CARRYB_27__2_), .CI(SUMB_27__3_), .CO(
        CARRYB_28__2_), .S(SUMB_28__2_) );
  ADDFX2 S2_28_1 ( .A(ab_28__1_), .B(CARRYB_27__1_), .CI(SUMB_27__2_), .CO(
        CARRYB_28__1_), .S(SUMB_28__1_) );
  ADDFX2 S2_27_3 ( .A(ab_27__3_), .B(CARRYB_26__3_), .CI(SUMB_26__4_), .CO(
        CARRYB_27__3_), .S(SUMB_27__3_) );
  ADDFX2 S2_27_2 ( .A(ab_27__2_), .B(CARRYB_26__2_), .CI(SUMB_26__3_), .CO(
        CARRYB_27__2_), .S(SUMB_27__2_) );
  ADDFX2 S2_27_1 ( .A(ab_27__1_), .B(CARRYB_26__1_), .CI(SUMB_26__2_), .CO(
        CARRYB_27__1_), .S(SUMB_27__1_) );
  ADDFX2 S1_25_0 ( .A(ab_25__0_), .B(CARRYB_24__0_), .CI(SUMB_24__1_), .CO(
        CARRYB_25__0_), .S(PRODUCT[25]) );
  ADDFX2 S2_26_4 ( .A(ab_26__4_), .B(CARRYB_25__4_), .CI(SUMB_25__5_), .CO(
        CARRYB_26__4_), .S(SUMB_26__4_) );
  ADDFX2 S2_26_3 ( .A(ab_26__3_), .B(CARRYB_25__3_), .CI(SUMB_25__4_), .CO(
        CARRYB_26__3_), .S(SUMB_26__3_) );
  ADDFX2 S2_26_2 ( .A(ab_26__2_), .B(CARRYB_25__2_), .CI(SUMB_25__3_), .CO(
        CARRYB_26__2_), .S(SUMB_26__2_) );
  ADDFX2 S2_26_1 ( .A(ab_26__1_), .B(CARRYB_25__1_), .CI(SUMB_25__2_), .CO(
        CARRYB_26__1_), .S(SUMB_26__1_) );
  ADDFX2 S1_24_0 ( .A(ab_24__0_), .B(CARRYB_23__0_), .CI(SUMB_23__1_), .CO(
        CARRYB_24__0_), .S(PRODUCT[24]) );
  ADDFX2 S2_25_5 ( .A(ab_25__5_), .B(CARRYB_24__5_), .CI(SUMB_24__6_), .CO(
        CARRYB_25__5_), .S(SUMB_25__5_) );
  ADDFX2 S2_25_4 ( .A(ab_25__4_), .B(CARRYB_24__4_), .CI(SUMB_24__5_), .CO(
        CARRYB_25__4_), .S(SUMB_25__4_) );
  ADDFX2 S2_25_3 ( .A(ab_25__3_), .B(CARRYB_24__3_), .CI(SUMB_24__4_), .CO(
        CARRYB_25__3_), .S(SUMB_25__3_) );
  ADDFX2 S2_25_2 ( .A(ab_25__2_), .B(CARRYB_24__2_), .CI(SUMB_24__3_), .CO(
        CARRYB_25__2_), .S(SUMB_25__2_) );
  ADDFX2 S2_25_1 ( .A(ab_25__1_), .B(CARRYB_24__1_), .CI(SUMB_24__2_), .CO(
        CARRYB_25__1_), .S(SUMB_25__1_) );
  ADDFX2 S1_23_0 ( .A(ab_23__0_), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(PRODUCT[23]) );
  ADDFX2 S2_24_6 ( .A(ab_24__6_), .B(CARRYB_23__6_), .CI(SUMB_23__7_), .CO(
        CARRYB_24__6_), .S(SUMB_24__6_) );
  ADDFX2 S2_24_5 ( .A(ab_24__5_), .B(CARRYB_23__5_), .CI(SUMB_23__6_), .CO(
        CARRYB_24__5_), .S(SUMB_24__5_) );
  ADDFX2 S2_24_4 ( .A(ab_24__4_), .B(CARRYB_23__4_), .CI(SUMB_23__5_), .CO(
        CARRYB_24__4_), .S(SUMB_24__4_) );
  ADDFX2 S2_24_3 ( .A(ab_24__3_), .B(CARRYB_23__3_), .CI(SUMB_23__4_), .CO(
        CARRYB_24__3_), .S(SUMB_24__3_) );
  ADDFX2 S2_24_2 ( .A(ab_24__2_), .B(CARRYB_23__2_), .CI(SUMB_23__3_), .CO(
        CARRYB_24__2_), .S(SUMB_24__2_) );
  ADDFX2 S2_24_1 ( .A(ab_24__1_), .B(CARRYB_23__1_), .CI(SUMB_23__2_), .CO(
        CARRYB_24__1_), .S(SUMB_24__1_) );
  ADDFX2 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(PRODUCT[22]) );
  ADDFX2 S2_23_6 ( .A(ab_23__6_), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  ADDFX2 S2_23_5 ( .A(ab_23__5_), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  ADDFX2 S2_23_4 ( .A(ab_23__4_), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  ADDFX2 S2_23_3 ( .A(ab_23__3_), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  ADDFX2 S2_23_2 ( .A(ab_23__2_), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  ADDFX2 S2_23_1 ( .A(ab_23__1_), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  ADDFX2 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(PRODUCT[21]) );
  ADDFX2 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  ADDFX2 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  ADDFX2 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  ADDFX2 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  ADDFX2 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  ADDFX2 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  ADDFX2 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(PRODUCT[20]) );
  ADDFX2 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  ADDFX2 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  ADDFX2 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  ADDFX2 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  ADDFX2 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  ADDFX2 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  ADDFX2 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(PRODUCT[19]) );
  ADDFX2 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  ADDFX2 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  ADDFX2 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  ADDFX2 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  ADDFX2 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  ADDFX2 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  ADDFX2 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  ADDFX2 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  ADDFX2 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  ADDFX2 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  ADDFX2 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  ADDFX2 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  ADDFX2 S2_6_6 ( .A(B[6]), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  ADDFX2 S2_5_5 ( .A(B[5]), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  XOR3X2 S2_29_2 ( .A(ab_29__2_), .B(CARRYB_28__2_), .C(SUMB_28__3_), .Y(
        SUMB_29__2_) );
  XOR3X2 S2_30_1 ( .A(ab_30__1_), .B(CARRYB_29__1_), .C(SUMB_29__2_), .Y(
        SUMB_30__1_) );
  ADDFX2 S2_2_13 ( .A(ab_2__13_), .B(n20), .CI(SUMB_1__14_), .CO(CARRYB_2__13_), .S(SUMB_2__13_) );
  ADDFX2 S2_2_11 ( .A(ab_2__11_), .B(n22), .CI(SUMB_1__12_), .CO(CARRYB_2__11_), .S(SUMB_2__11_) );
  ADDFX2 S2_2_15 ( .A(ab_2__15_), .B(n18), .CI(SUMB_1__16_), .CO(CARRYB_2__15_), .S(SUMB_2__15_) );
  ADDFX2 S2_2_14 ( .A(ab_2__14_), .B(n21), .CI(SUMB_1__15_), .CO(CARRYB_2__14_), .S(SUMB_2__14_) );
  ADDFX2 S2_2_12 ( .A(ab_2__12_), .B(n19), .CI(SUMB_1__13_), .CO(CARRYB_2__12_), .S(SUMB_2__12_) );
  ADDFX2 S2_2_10 ( .A(ab_2__10_), .B(n14), .CI(SUMB_1__11_), .CO(CARRYB_2__10_), .S(SUMB_2__10_) );
  ADDFX2 S2_2_9 ( .A(ab_2__9_), .B(n13), .CI(SUMB_1__10_), .CO(CARRYB_2__9_), 
        .S(SUMB_2__9_) );
  ADDFX2 S2_2_8 ( .A(ab_2__8_), .B(n17), .CI(SUMB_1__9_), .CO(CARRYB_2__8_), 
        .S(SUMB_2__8_) );
  ADDFX2 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), 
        .CO(CARRYB_14__13_), .S(SUMB_14__13_) );
  ADDFX2 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), 
        .CO(CARRYB_14__12_), .S(SUMB_14__12_) );
  ADDFX2 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), 
        .CO(CARRYB_14__11_), .S(SUMB_14__11_) );
  ADDFX2 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  ADDFX2 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  ADDFX2 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), 
        .CO(CARRYB_15__14_), .S(SUMB_15__14_) );
  ADDFX2 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), 
        .CO(CARRYB_15__13_), .S(SUMB_15__13_) );
  ADDFX2 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), 
        .CO(CARRYB_15__12_), .S(SUMB_15__12_) );
  ADDFX2 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), 
        .CO(CARRYB_14__15_), .S(SUMB_14__15_) );
  ADDFX2 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), 
        .CO(CARRYB_15__11_), .S(SUMB_15__11_) );
  ADDFX2 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), 
        .CO(CARRYB_15__10_), .S(SUMB_15__10_) );
  ADDFX2 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  ADDFX2 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  ADDFX2 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  ADDFX2 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), 
        .CO(CARRYB_14__10_), .S(SUMB_14__10_) );
  ADDFX2 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  ADDFX2 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  ADDFX2 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  ADDFX2 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), 
        .CO(CARRYB_13__15_), .S(SUMB_13__15_) );
  ADDFX2 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), 
        .CO(CARRYB_13__14_), .S(SUMB_13__14_) );
  ADDFX2 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), 
        .CO(CARRYB_13__12_), .S(SUMB_13__12_) );
  ADDFX2 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), 
        .CO(CARRYB_13__11_), .S(SUMB_13__11_) );
  ADDFX2 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), 
        .CO(CARRYB_13__10_), .S(SUMB_13__10_) );
  ADDFX2 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  ADDFX2 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  ADDFX2 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  ADDFX2 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), 
        .CO(CARRYB_12__15_), .S(SUMB_12__15_) );
  ADDFX2 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), 
        .CO(CARRYB_12__14_), .S(SUMB_12__14_) );
  ADDFX2 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), 
        .CO(CARRYB_12__13_), .S(SUMB_12__13_) );
  ADDFX2 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), 
        .CO(CARRYB_12__11_), .S(SUMB_12__11_) );
  ADDFX2 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), 
        .CO(CARRYB_12__10_), .S(SUMB_12__10_) );
  ADDFX2 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  ADDFX2 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), 
        .CO(CARRYB_11__15_), .S(SUMB_11__15_) );
  ADDFX2 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), 
        .CO(CARRYB_11__14_), .S(SUMB_11__14_) );
  ADDFX2 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), 
        .CO(CARRYB_11__13_), .S(SUMB_11__13_) );
  ADDFX2 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), 
        .CO(CARRYB_11__12_), .S(SUMB_11__12_) );
  ADDFX2 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), 
        .CO(CARRYB_11__10_), .S(SUMB_11__10_) );
  ADDFX2 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  ADDFX2 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  ADDFX2 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  ADDFX2 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  ADDFX2 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  ADDFX2 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  ADDFX2 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  ADDFX2 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  ADDFX2 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  ADDFX2 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  ADDFX2 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  ADDFX2 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  ADDFX2 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  ADDFX2 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  ADDFX2 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  ADDFX2 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  ADDFX2 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  ADDFX2 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  ADDFX2 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  ADDFX2 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  ADDFX2 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  ADDFX2 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  ADDFX2 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  ADDFX2 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  ADDFX2 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  ADDFX2 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  ADDFX2 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  ADDFX2 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  ADDFX2 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  ADDFX2 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  ADDFX2 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  ADDFX2 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  ADDFX2 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  ADDFX2 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  ADDFX2 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  ADDFX2 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  ADDFX2 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  ADDFX2 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  ADDFX2 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  ADDFX2 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  ADDFX2 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  ADDFX2 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  ADDFX2 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  ADDFX2 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  ADDFX2 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  ADDFX2 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  ADDFX2 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  ADDFX2 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  ADDFX2 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  ADDFX2 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  ADDFX2 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  ADDFX2 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  ADDFX2 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  ADDFX2 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  ADDFX2 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  ADDFX2 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  ADDFX2 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  ADDFX2 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  ADDFX2 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  ADDFX2 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  ADDFX2 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  ADDFX2 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  ADDFX2 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  ADDFX2 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  ADDFX2 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  ADDFX2 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  ADDFX2 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  ADDFX2 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  ADDFX2 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  ADDFX2 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  ADDFX2 S2_2_7 ( .A(ab_2__7_), .B(n16), .CI(SUMB_1__8_), .CO(CARRYB_2__7_), 
        .S(SUMB_2__7_) );
  ADDFX2 S2_2_6 ( .A(ab_2__6_), .B(n15), .CI(SUMB_1__7_), .CO(CARRYB_2__6_), 
        .S(SUMB_2__6_) );
  ADDFX2 S2_2_5 ( .A(ab_2__5_), .B(n9), .CI(SUMB_1__6_), .CO(CARRYB_2__5_), 
        .S(SUMB_2__5_) );
  ADDFX2 S1_2_0 ( .A(ab_2__0_), .B(n7), .CI(SUMB_1__1_), .CO(CARRYB_2__0_), 
        .S(PRODUCT[2]) );
  ADDFX2 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(PRODUCT[3]) );
  ADDFX2 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(PRODUCT[4]) );
  ADDFX2 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(PRODUCT[5]) );
  ADDFX2 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(PRODUCT[15]) );
  ADDFX2 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(PRODUCT[14]) );
  ADDFX2 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  ADDFX2 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  ADDFX2 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  ADDFX2 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  ADDFX2 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  ADDFX2 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  ADDFX2 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(PRODUCT[13]) );
  ADDFX2 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  ADDFX2 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  ADDFX2 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  ADDFX2 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  ADDFX2 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  ADDFX2 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  ADDFX2 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(PRODUCT[12]) );
  ADDFX2 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  ADDFX2 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  ADDFX2 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  ADDFX2 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  ADDFX2 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  ADDFX2 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  ADDFX2 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(PRODUCT[11]) );
  ADDFX2 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  ADDFX2 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  ADDFX2 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  ADDFX2 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  ADDFX2 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  ADDFX2 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  ADDFX2 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(PRODUCT[10]) );
  ADDFX2 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  ADDFX2 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  ADDFX2 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  ADDFX2 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  ADDFX2 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  ADDFX2 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  ADDFX2 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(PRODUCT[9]) );
  ADDFX2 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  ADDFX2 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  ADDFX2 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  ADDFX2 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  ADDFX2 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  ADDFX2 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  ADDFX2 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(PRODUCT[8]) );
  ADDFX2 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  ADDFX2 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  ADDFX2 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  ADDFX2 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  ADDFX2 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  ADDFX2 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  ADDFX2 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(PRODUCT[7]) );
  ADDFX2 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  ADDFX2 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  ADDFX2 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  ADDFX2 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  ADDFX2 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  ADDFX2 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  ADDFX2 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(PRODUCT[6]) );
  ADDFX2 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  ADDFX2 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  ADDFX2 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  ADDFX2 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  ADDFX2 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  ADDFX2 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  ADDFX2 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  ADDFX2 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  ADDFX2 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  ADDFX2 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  ADDFX2 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  ADDFX2 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  ADDFX2 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  ADDFX2 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  ADDFX2 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  ADDFX2 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  ADDFX2 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  ADDFX2 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  ADDFX2 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  ADDFX2 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  ADDFX2 S2_2_4 ( .A(ab_2__4_), .B(n8), .CI(SUMB_1__5_), .CO(CARRYB_2__4_), 
        .S(SUMB_2__4_) );
  ADDFX2 S2_2_3 ( .A(ab_2__3_), .B(n12), .CI(SUMB_1__4_), .CO(CARRYB_2__3_), 
        .S(SUMB_2__3_) );
  ADDFX2 S2_2_2 ( .A(n44), .B(n11), .CI(SUMB_1__3_), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  ADDFX2 S2_2_1 ( .A(ab_2__1_), .B(n10), .CI(SUMB_1__2_), .CO(CARRYB_2__1_), 
        .S(SUMB_2__1_) );
  ADDFX2 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  ADDFX2 S2_4_4 ( .A(n52), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(CARRYB_4__4_), .S(SUMB_4__4_) );
  ADDFX2 S2_3_3 ( .A(n48), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(CARRYB_3__3_), .S(SUMB_3__3_) );
  ADDFX2 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  ADDFX2 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  ADDFX2 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  ADDFX2 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  ADDFX2 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  AND2X2 U2 ( .A(ab_0__1_), .B(ab_1__0_), .Y(n7) );
  AND2X2 U3 ( .A(ab_0__5_), .B(ab_1__4_), .Y(n8) );
  AND2X2 U4 ( .A(ab_0__6_), .B(ab_1__5_), .Y(n9) );
  AND2X2 U5 ( .A(ab_0__2_), .B(n40), .Y(n10) );
  AND2X2 U6 ( .A(ab_0__3_), .B(ab_1__2_), .Y(n11) );
  AND2X2 U7 ( .A(ab_0__4_), .B(ab_1__3_), .Y(n12) );
  AND2X2 U8 ( .A(ab_0__10_), .B(ab_1__9_), .Y(n13) );
  AND2X2 U9 ( .A(ab_0__11_), .B(ab_1__10_), .Y(n14) );
  AND2X2 U10 ( .A(ab_0__7_), .B(ab_1__6_), .Y(n15) );
  AND2X2 U11 ( .A(ab_0__8_), .B(ab_1__7_), .Y(n16) );
  AND2X2 U12 ( .A(ab_0__9_), .B(ab_1__8_), .Y(n17) );
  AND2X2 U13 ( .A(ab_0__16_), .B(ab_1__15_), .Y(n18) );
  AND2X2 U14 ( .A(ab_0__13_), .B(ab_1__12_), .Y(n19) );
  AND2X2 U15 ( .A(ab_0__14_), .B(ab_1__13_), .Y(n20) );
  AND2X2 U16 ( .A(ab_0__15_), .B(ab_1__14_), .Y(n21) );
  AND2X2 U17 ( .A(ab_0__12_), .B(ab_1__11_), .Y(n22) );
  AND2X2 U18 ( .A(ab_0__17_), .B(ab_1__16_), .Y(n23) );
  AND2X2 U19 ( .A(ab_0__18_), .B(ab_1__17_), .Y(n24) );
  AND2X2 U20 ( .A(ab_0__19_), .B(ab_1__18_), .Y(n25) );
  AND2X2 U21 ( .A(ab_0__20_), .B(ab_1__19_), .Y(n26) );
  AND2X2 U22 ( .A(ab_0__21_), .B(ab_1__20_), .Y(n27) );
  AND2X2 U23 ( .A(ab_0__22_), .B(ab_1__21_), .Y(n28) );
  AND2X2 U24 ( .A(ab_0__23_), .B(ab_1__22_), .Y(n29) );
  AND2X2 U25 ( .A(ab_0__24_), .B(ab_1__23_), .Y(n30) );
  AND2X2 U26 ( .A(ab_0__25_), .B(ab_1__24_), .Y(n31) );
  AND2X2 U27 ( .A(ab_0__26_), .B(ab_1__25_), .Y(n32) );
  AND2X2 U28 ( .A(ab_0__27_), .B(ab_1__26_), .Y(n33) );
  AND2X2 U29 ( .A(ab_0__28_), .B(ab_1__27_), .Y(n34) );
  AND2X2 U30 ( .A(ab_0__29_), .B(ab_1__28_), .Y(n35) );
  AND2X2 U31 ( .A(ab_0__30_), .B(ab_1__29_), .Y(n36) );
  XOR2X1 U32 ( .A(ab_1__2_), .B(ab_0__3_), .Y(SUMB_1__2_) );
  XOR2X1 U33 ( .A(ab_1__3_), .B(ab_0__4_), .Y(SUMB_1__3_) );
  XOR2X1 U34 ( .A(ab_1__4_), .B(ab_0__5_), .Y(SUMB_1__4_) );
  XOR2X1 U35 ( .A(ab_1__5_), .B(ab_0__6_), .Y(SUMB_1__5_) );
  INVX1 U36 ( .A(n44), .Y(n45) );
  INVX1 U37 ( .A(n48), .Y(n49) );
  INVX1 U38 ( .A(n52), .Y(n54) );
  INVX1 U39 ( .A(A[3]), .Y(n51) );
  INVX1 U40 ( .A(A[4]), .Y(n55) );
  INVX1 U41 ( .A(A[1]), .Y(n43) );
  INVX1 U42 ( .A(A[2]), .Y(n47) );
  INVX1 U43 ( .A(n44), .Y(n46) );
  INVX1 U44 ( .A(n48), .Y(n50) );
  INVX1 U45 ( .A(A[1]), .Y(n42) );
  INVX1 U46 ( .A(n40), .Y(n41) );
  XOR2X1 U47 ( .A(n40), .B(ab_0__2_), .Y(SUMB_1__1_) );
  XOR2X1 U48 ( .A(ab_1__6_), .B(ab_0__7_), .Y(SUMB_1__6_) );
  XOR2X1 U49 ( .A(ab_1__7_), .B(ab_0__8_), .Y(SUMB_1__7_) );
  XOR2X1 U50 ( .A(ab_1__8_), .B(ab_0__9_), .Y(SUMB_1__8_) );
  INVX1 U51 ( .A(n47), .Y(n44) );
  INVX1 U52 ( .A(n51), .Y(n48) );
  INVX1 U53 ( .A(n53), .Y(n52) );
  XOR2X1 U54 ( .A(ab_1__9_), .B(ab_0__10_), .Y(SUMB_1__9_) );
  XOR2X1 U55 ( .A(ab_1__10_), .B(ab_0__11_), .Y(SUMB_1__10_) );
  XOR2X1 U56 ( .A(ab_1__11_), .B(ab_0__12_), .Y(SUMB_1__11_) );
  XOR2X1 U57 ( .A(ab_1__13_), .B(ab_0__14_), .Y(SUMB_1__13_) );
  XOR2X1 U58 ( .A(ab_1__15_), .B(ab_0__16_), .Y(SUMB_1__15_) );
  XOR2X1 U59 ( .A(ab_1__16_), .B(ab_0__17_), .Y(SUMB_1__16_) );
  XOR2X1 U60 ( .A(ab_1__12_), .B(ab_0__13_), .Y(SUMB_1__12_) );
  XOR2X1 U61 ( .A(ab_1__14_), .B(ab_0__15_), .Y(SUMB_1__14_) );
  INVX1 U62 ( .A(n43), .Y(n40) );
  XOR2X1 U63 ( .A(CARRYB_30__0_), .B(SUMB_30__1_), .Y(PRODUCT[31]) );
  INVX1 U64 ( .A(B[4]), .Y(n53) );
  XOR2X1 U65 ( .A(ab_1__17_), .B(ab_0__18_), .Y(SUMB_1__17_) );
  XOR2X1 U66 ( .A(ab_1__18_), .B(ab_0__19_), .Y(SUMB_1__18_) );
  XOR2X1 U67 ( .A(ab_1__19_), .B(ab_0__20_), .Y(SUMB_1__19_) );
  XOR2X1 U68 ( .A(ab_1__20_), .B(ab_0__21_), .Y(SUMB_1__20_) );
  XOR2X1 U69 ( .A(ab_1__21_), .B(ab_0__22_), .Y(SUMB_1__21_) );
  XOR2X1 U70 ( .A(ab_1__22_), .B(ab_0__23_), .Y(SUMB_1__22_) );
  XOR2X1 U71 ( .A(ab_1__23_), .B(ab_0__24_), .Y(SUMB_1__23_) );
  XOR2X1 U72 ( .A(ab_1__24_), .B(ab_0__25_), .Y(SUMB_1__24_) );
  XOR2X1 U73 ( .A(ab_1__25_), .B(ab_0__26_), .Y(SUMB_1__25_) );
  XOR2X1 U74 ( .A(ab_1__26_), .B(ab_0__27_), .Y(SUMB_1__26_) );
  XOR2X1 U75 ( .A(ab_1__27_), .B(ab_0__28_), .Y(SUMB_1__27_) );
  XOR2X1 U76 ( .A(ab_1__28_), .B(ab_0__29_), .Y(SUMB_1__28_) );
  XOR2X1 U77 ( .A(ab_1__29_), .B(ab_0__30_), .Y(SUMB_1__29_) );
  INVX1 U78 ( .A(B[7]), .Y(n58) );
  INVX1 U79 ( .A(B[0]), .Y(n38) );
  INVX1 U80 ( .A(B[11]), .Y(n63) );
  INVX1 U81 ( .A(B[0]), .Y(n37) );
  INVX1 U82 ( .A(B[8]), .Y(n59) );
  INVX1 U83 ( .A(B[9]), .Y(n60) );
  INVX1 U84 ( .A(B[10]), .Y(n62) );
  INVX1 U85 ( .A(B[13]), .Y(n65) );
  INVX1 U86 ( .A(B[15]), .Y(n67) );
  INVX1 U87 ( .A(B[14]), .Y(n66) );
  INVX1 U88 ( .A(B[0]), .Y(n39) );
  INVX1 U89 ( .A(B[9]), .Y(n61) );
  INVX1 U90 ( .A(B[5]), .Y(n56) );
  INVX1 U91 ( .A(B[6]), .Y(n57) );
  INVX1 U92 ( .A(B[12]), .Y(n64) );
  XOR2X1 U93 ( .A(ab_1__0_), .B(ab_0__1_), .Y(PRODUCT[1]) );
  INVX1 U94 ( .A(B[16]), .Y(n69) );
  INVX1 U95 ( .A(B[17]), .Y(n70) );
  INVX1 U96 ( .A(B[18]), .Y(n71) );
  INVX1 U97 ( .A(B[19]), .Y(n72) );
  INVX1 U98 ( .A(B[20]), .Y(n73) );
  INVX1 U99 ( .A(B[21]), .Y(n74) );
  INVX1 U100 ( .A(B[22]), .Y(n75) );
  INVX1 U101 ( .A(B[23]), .Y(n76) );
  INVX1 U102 ( .A(B[24]), .Y(n77) );
  INVX1 U103 ( .A(B[25]), .Y(n78) );
  INVX1 U104 ( .A(B[26]), .Y(n79) );
  INVX1 U105 ( .A(B[27]), .Y(n80) );
  INVX1 U106 ( .A(B[28]), .Y(n81) );
  INVX1 U107 ( .A(B[29]), .Y(n82) );
  INVX1 U108 ( .A(B[30]), .Y(n68) );
  NOR2X1 U109 ( .A(n60), .B(n59), .Y(ab_9__8_) );
  NOR2X1 U110 ( .A(n61), .B(n58), .Y(ab_9__7_) );
  NOR2X1 U111 ( .A(n60), .B(n57), .Y(ab_9__6_) );
  NOR2X1 U112 ( .A(n60), .B(n56), .Y(ab_9__5_) );
  NOR2X1 U113 ( .A(n60), .B(n55), .Y(ab_9__4_) );
  NOR2X1 U114 ( .A(n60), .B(n51), .Y(ab_9__3_) );
  NOR2X1 U115 ( .A(n60), .B(n47), .Y(ab_9__2_) );
  NOR2X1 U116 ( .A(n60), .B(n75), .Y(ab_9__22_) );
  NOR2X1 U117 ( .A(n61), .B(n74), .Y(ab_9__21_) );
  NOR2X1 U118 ( .A(n61), .B(n73), .Y(ab_9__20_) );
  NOR2X1 U119 ( .A(n60), .B(n43), .Y(ab_9__1_) );
  NOR2X1 U120 ( .A(n60), .B(n72), .Y(ab_9__19_) );
  NOR2X1 U121 ( .A(n61), .B(n71), .Y(ab_9__18_) );
  NOR2X1 U122 ( .A(n60), .B(n70), .Y(ab_9__17_) );
  NOR2X1 U123 ( .A(n61), .B(n69), .Y(ab_9__16_) );
  NOR2X1 U124 ( .A(n60), .B(n67), .Y(ab_9__15_) );
  NOR2X1 U125 ( .A(n61), .B(n66), .Y(ab_9__14_) );
  NOR2X1 U126 ( .A(n60), .B(n65), .Y(ab_9__13_) );
  NOR2X1 U127 ( .A(n61), .B(n64), .Y(ab_9__12_) );
  NOR2X1 U128 ( .A(n60), .B(n63), .Y(ab_9__11_) );
  NOR2X1 U129 ( .A(n61), .B(n62), .Y(ab_9__10_) );
  NOR2X1 U130 ( .A(n60), .B(n37), .Y(ab_9__0_) );
  NOR2X1 U131 ( .A(n60), .B(n59), .Y(ab_8__9_) );
  NOR2X1 U132 ( .A(n58), .B(n59), .Y(ab_8__7_) );
  NOR2X1 U133 ( .A(n57), .B(n59), .Y(ab_8__6_) );
  NOR2X1 U134 ( .A(n56), .B(n59), .Y(ab_8__5_) );
  NOR2X1 U135 ( .A(n55), .B(n59), .Y(ab_8__4_) );
  NOR2X1 U136 ( .A(n51), .B(n59), .Y(ab_8__3_) );
  NOR2X1 U137 ( .A(n47), .B(n59), .Y(ab_8__2_) );
  NOR2X1 U138 ( .A(n76), .B(n59), .Y(ab_8__23_) );
  NOR2X1 U139 ( .A(n75), .B(n59), .Y(ab_8__22_) );
  NOR2X1 U140 ( .A(n74), .B(n59), .Y(ab_8__21_) );
  NOR2X1 U141 ( .A(n73), .B(n59), .Y(ab_8__20_) );
  NOR2X1 U142 ( .A(n43), .B(n59), .Y(ab_8__1_) );
  NOR2X1 U143 ( .A(n72), .B(n59), .Y(ab_8__19_) );
  NOR2X1 U144 ( .A(n71), .B(n59), .Y(ab_8__18_) );
  NOR2X1 U145 ( .A(n70), .B(n59), .Y(ab_8__17_) );
  NOR2X1 U146 ( .A(n69), .B(n59), .Y(ab_8__16_) );
  NOR2X1 U147 ( .A(n67), .B(n59), .Y(ab_8__15_) );
  NOR2X1 U148 ( .A(n66), .B(n59), .Y(ab_8__14_) );
  NOR2X1 U149 ( .A(n65), .B(n59), .Y(ab_8__13_) );
  NOR2X1 U150 ( .A(n64), .B(n59), .Y(ab_8__12_) );
  NOR2X1 U151 ( .A(n63), .B(n59), .Y(ab_8__11_) );
  NOR2X1 U152 ( .A(n62), .B(n59), .Y(ab_8__10_) );
  NOR2X1 U153 ( .A(n39), .B(n59), .Y(ab_8__0_) );
  NOR2X1 U154 ( .A(n60), .B(n58), .Y(ab_7__9_) );
  NOR2X1 U155 ( .A(n59), .B(n58), .Y(ab_7__8_) );
  NOR2X1 U156 ( .A(n57), .B(n58), .Y(ab_7__6_) );
  NOR2X1 U157 ( .A(n56), .B(n58), .Y(ab_7__5_) );
  NOR2X1 U158 ( .A(n55), .B(n58), .Y(ab_7__4_) );
  NOR2X1 U159 ( .A(n51), .B(n58), .Y(ab_7__3_) );
  NOR2X1 U160 ( .A(n47), .B(n58), .Y(ab_7__2_) );
  NOR2X1 U161 ( .A(n77), .B(n58), .Y(ab_7__24_) );
  NOR2X1 U162 ( .A(n76), .B(n58), .Y(ab_7__23_) );
  NOR2X1 U163 ( .A(n75), .B(n58), .Y(ab_7__22_) );
  NOR2X1 U164 ( .A(n74), .B(n58), .Y(ab_7__21_) );
  NOR2X1 U165 ( .A(n73), .B(n58), .Y(ab_7__20_) );
  NOR2X1 U166 ( .A(n43), .B(n58), .Y(ab_7__1_) );
  NOR2X1 U167 ( .A(n72), .B(n58), .Y(ab_7__19_) );
  NOR2X1 U168 ( .A(n71), .B(n58), .Y(ab_7__18_) );
  NOR2X1 U169 ( .A(n70), .B(n58), .Y(ab_7__17_) );
  NOR2X1 U170 ( .A(n69), .B(n58), .Y(ab_7__16_) );
  NOR2X1 U171 ( .A(n67), .B(n58), .Y(ab_7__15_) );
  NOR2X1 U172 ( .A(n66), .B(n58), .Y(ab_7__14_) );
  NOR2X1 U173 ( .A(n65), .B(n58), .Y(ab_7__13_) );
  NOR2X1 U174 ( .A(n64), .B(n58), .Y(ab_7__12_) );
  NOR2X1 U175 ( .A(n63), .B(n58), .Y(ab_7__11_) );
  NOR2X1 U176 ( .A(n62), .B(n58), .Y(ab_7__10_) );
  NOR2X1 U177 ( .A(n37), .B(n58), .Y(ab_7__0_) );
  NOR2X1 U178 ( .A(n60), .B(n57), .Y(ab_6__9_) );
  NOR2X1 U179 ( .A(n59), .B(n57), .Y(ab_6__8_) );
  NOR2X1 U180 ( .A(n58), .B(n57), .Y(ab_6__7_) );
  NOR2X1 U181 ( .A(n56), .B(n57), .Y(ab_6__5_) );
  NOR2X1 U182 ( .A(n55), .B(n57), .Y(ab_6__4_) );
  NOR2X1 U183 ( .A(n51), .B(n57), .Y(ab_6__3_) );
  NOR2X1 U184 ( .A(n47), .B(n57), .Y(ab_6__2_) );
  NOR2X1 U185 ( .A(n78), .B(n57), .Y(ab_6__25_) );
  NOR2X1 U186 ( .A(n77), .B(n57), .Y(ab_6__24_) );
  NOR2X1 U187 ( .A(n76), .B(n57), .Y(ab_6__23_) );
  NOR2X1 U188 ( .A(n75), .B(n57), .Y(ab_6__22_) );
  NOR2X1 U189 ( .A(n74), .B(n57), .Y(ab_6__21_) );
  NOR2X1 U190 ( .A(n73), .B(n57), .Y(ab_6__20_) );
  NOR2X1 U191 ( .A(n43), .B(n57), .Y(ab_6__1_) );
  NOR2X1 U192 ( .A(n72), .B(n57), .Y(ab_6__19_) );
  NOR2X1 U193 ( .A(n71), .B(n57), .Y(ab_6__18_) );
  NOR2X1 U194 ( .A(n70), .B(n57), .Y(ab_6__17_) );
  NOR2X1 U195 ( .A(n69), .B(n57), .Y(ab_6__16_) );
  NOR2X1 U196 ( .A(n67), .B(n57), .Y(ab_6__15_) );
  NOR2X1 U197 ( .A(n66), .B(n57), .Y(ab_6__14_) );
  NOR2X1 U198 ( .A(n65), .B(n57), .Y(ab_6__13_) );
  NOR2X1 U199 ( .A(n64), .B(n57), .Y(ab_6__12_) );
  NOR2X1 U200 ( .A(n63), .B(n57), .Y(ab_6__11_) );
  NOR2X1 U201 ( .A(n62), .B(n57), .Y(ab_6__10_) );
  NOR2X1 U202 ( .A(n37), .B(n57), .Y(ab_6__0_) );
  NOR2X1 U203 ( .A(n60), .B(n56), .Y(ab_5__9_) );
  NOR2X1 U204 ( .A(n59), .B(n56), .Y(ab_5__8_) );
  NOR2X1 U205 ( .A(n58), .B(n56), .Y(ab_5__7_) );
  NOR2X1 U206 ( .A(n57), .B(n56), .Y(ab_5__6_) );
  NOR2X1 U207 ( .A(n55), .B(n56), .Y(ab_5__4_) );
  NOR2X1 U208 ( .A(n50), .B(n56), .Y(ab_5__3_) );
  NOR2X1 U209 ( .A(n47), .B(n56), .Y(ab_5__2_) );
  NOR2X1 U210 ( .A(n79), .B(n56), .Y(ab_5__26_) );
  NOR2X1 U211 ( .A(n78), .B(n56), .Y(ab_5__25_) );
  NOR2X1 U212 ( .A(n77), .B(n56), .Y(ab_5__24_) );
  NOR2X1 U213 ( .A(n76), .B(n56), .Y(ab_5__23_) );
  NOR2X1 U214 ( .A(n75), .B(n56), .Y(ab_5__22_) );
  NOR2X1 U215 ( .A(n74), .B(n56), .Y(ab_5__21_) );
  NOR2X1 U216 ( .A(n73), .B(n56), .Y(ab_5__20_) );
  NOR2X1 U217 ( .A(n43), .B(n56), .Y(ab_5__1_) );
  NOR2X1 U218 ( .A(n72), .B(n56), .Y(ab_5__19_) );
  NOR2X1 U219 ( .A(n71), .B(n56), .Y(ab_5__18_) );
  NOR2X1 U220 ( .A(n70), .B(n56), .Y(ab_5__17_) );
  NOR2X1 U221 ( .A(n69), .B(n56), .Y(ab_5__16_) );
  NOR2X1 U222 ( .A(n67), .B(n56), .Y(ab_5__15_) );
  NOR2X1 U223 ( .A(n66), .B(n56), .Y(ab_5__14_) );
  NOR2X1 U224 ( .A(n65), .B(n56), .Y(ab_5__13_) );
  NOR2X1 U225 ( .A(n64), .B(n56), .Y(ab_5__12_) );
  NOR2X1 U226 ( .A(n63), .B(n56), .Y(ab_5__11_) );
  NOR2X1 U227 ( .A(n62), .B(n56), .Y(ab_5__10_) );
  NOR2X1 U228 ( .A(n37), .B(n56), .Y(ab_5__0_) );
  NOR2X1 U229 ( .A(n60), .B(n55), .Y(ab_4__9_) );
  NOR2X1 U230 ( .A(n59), .B(n55), .Y(ab_4__8_) );
  NOR2X1 U231 ( .A(n58), .B(n55), .Y(ab_4__7_) );
  NOR2X1 U232 ( .A(n57), .B(n55), .Y(ab_4__6_) );
  NOR2X1 U233 ( .A(n56), .B(n55), .Y(ab_4__5_) );
  NOR2X1 U234 ( .A(n50), .B(n55), .Y(ab_4__3_) );
  NOR2X1 U235 ( .A(n46), .B(n55), .Y(ab_4__2_) );
  NOR2X1 U236 ( .A(n80), .B(n55), .Y(ab_4__27_) );
  NOR2X1 U237 ( .A(n79), .B(n55), .Y(ab_4__26_) );
  NOR2X1 U238 ( .A(n78), .B(n55), .Y(ab_4__25_) );
  NOR2X1 U239 ( .A(n77), .B(n55), .Y(ab_4__24_) );
  NOR2X1 U240 ( .A(n76), .B(n55), .Y(ab_4__23_) );
  NOR2X1 U241 ( .A(n75), .B(n55), .Y(ab_4__22_) );
  NOR2X1 U242 ( .A(n74), .B(n55), .Y(ab_4__21_) );
  NOR2X1 U243 ( .A(n73), .B(n55), .Y(ab_4__20_) );
  NOR2X1 U244 ( .A(n43), .B(n55), .Y(ab_4__1_) );
  NOR2X1 U245 ( .A(n72), .B(n55), .Y(ab_4__19_) );
  NOR2X1 U246 ( .A(n71), .B(n55), .Y(ab_4__18_) );
  NOR2X1 U247 ( .A(n70), .B(n55), .Y(ab_4__17_) );
  NOR2X1 U248 ( .A(n69), .B(n55), .Y(ab_4__16_) );
  NOR2X1 U249 ( .A(n67), .B(n55), .Y(ab_4__15_) );
  NOR2X1 U250 ( .A(n66), .B(n55), .Y(ab_4__14_) );
  NOR2X1 U251 ( .A(n65), .B(n55), .Y(ab_4__13_) );
  NOR2X1 U252 ( .A(n64), .B(n55), .Y(ab_4__12_) );
  NOR2X1 U253 ( .A(n63), .B(n55), .Y(ab_4__11_) );
  NOR2X1 U254 ( .A(n62), .B(n55), .Y(ab_4__10_) );
  NOR2X1 U255 ( .A(n37), .B(n55), .Y(ab_4__0_) );
  NOR2X1 U256 ( .A(n60), .B(n50), .Y(ab_3__9_) );
  NOR2X1 U257 ( .A(n59), .B(n50), .Y(ab_3__8_) );
  NOR2X1 U258 ( .A(n58), .B(n50), .Y(ab_3__7_) );
  NOR2X1 U259 ( .A(n57), .B(n50), .Y(ab_3__6_) );
  NOR2X1 U260 ( .A(n56), .B(n50), .Y(ab_3__5_) );
  NOR2X1 U261 ( .A(n55), .B(n50), .Y(ab_3__4_) );
  NOR2X1 U262 ( .A(n46), .B(n50), .Y(ab_3__2_) );
  NOR2X1 U263 ( .A(n81), .B(n50), .Y(ab_3__28_) );
  NOR2X1 U264 ( .A(n80), .B(n50), .Y(ab_3__27_) );
  NOR2X1 U265 ( .A(n79), .B(n50), .Y(ab_3__26_) );
  NOR2X1 U266 ( .A(n78), .B(n50), .Y(ab_3__25_) );
  NOR2X1 U267 ( .A(n77), .B(n50), .Y(ab_3__24_) );
  NOR2X1 U268 ( .A(n76), .B(n50), .Y(ab_3__23_) );
  NOR2X1 U269 ( .A(n75), .B(n50), .Y(ab_3__22_) );
  NOR2X1 U270 ( .A(n74), .B(n50), .Y(ab_3__21_) );
  NOR2X1 U271 ( .A(n73), .B(n50), .Y(ab_3__20_) );
  NOR2X1 U272 ( .A(n42), .B(n50), .Y(ab_3__1_) );
  NOR2X1 U273 ( .A(n72), .B(n50), .Y(ab_3__19_) );
  NOR2X1 U274 ( .A(n71), .B(n51), .Y(ab_3__18_) );
  NOR2X1 U275 ( .A(n70), .B(n51), .Y(ab_3__17_) );
  NOR2X1 U276 ( .A(n69), .B(n51), .Y(ab_3__16_) );
  NOR2X1 U277 ( .A(n67), .B(n51), .Y(ab_3__15_) );
  NOR2X1 U278 ( .A(n66), .B(n51), .Y(ab_3__14_) );
  NOR2X1 U279 ( .A(n65), .B(n51), .Y(ab_3__13_) );
  NOR2X1 U280 ( .A(n64), .B(n51), .Y(ab_3__12_) );
  NOR2X1 U281 ( .A(n63), .B(n51), .Y(ab_3__11_) );
  NOR2X1 U282 ( .A(n62), .B(n51), .Y(ab_3__10_) );
  NOR2X1 U283 ( .A(n37), .B(n51), .Y(ab_3__0_) );
  NOR2X1 U284 ( .A(n42), .B(n68), .Y(ab_30__1_) );
  NOR2X1 U285 ( .A(n37), .B(n68), .Y(ab_30__0_) );
  NOR2X1 U286 ( .A(n60), .B(n46), .Y(ab_2__9_) );
  NOR2X1 U287 ( .A(n59), .B(n46), .Y(ab_2__8_) );
  NOR2X1 U288 ( .A(n58), .B(n46), .Y(ab_2__7_) );
  NOR2X1 U289 ( .A(n57), .B(n46), .Y(ab_2__6_) );
  NOR2X1 U290 ( .A(n56), .B(n46), .Y(ab_2__5_) );
  NOR2X1 U291 ( .A(n55), .B(n46), .Y(ab_2__4_) );
  NOR2X1 U292 ( .A(n50), .B(n46), .Y(ab_2__3_) );
  NOR2X1 U293 ( .A(n82), .B(n47), .Y(ab_2__29_) );
  NOR2X1 U294 ( .A(n81), .B(n47), .Y(ab_2__28_) );
  NOR2X1 U295 ( .A(n80), .B(n47), .Y(ab_2__27_) );
  NOR2X1 U296 ( .A(n79), .B(n45), .Y(ab_2__26_) );
  NOR2X1 U297 ( .A(n78), .B(n46), .Y(ab_2__25_) );
  NOR2X1 U298 ( .A(n77), .B(n46), .Y(ab_2__24_) );
  NOR2X1 U299 ( .A(n76), .B(n46), .Y(ab_2__23_) );
  NOR2X1 U300 ( .A(n75), .B(n46), .Y(ab_2__22_) );
  NOR2X1 U301 ( .A(n74), .B(n46), .Y(ab_2__21_) );
  NOR2X1 U302 ( .A(n73), .B(n46), .Y(ab_2__20_) );
  NOR2X1 U303 ( .A(n42), .B(n46), .Y(ab_2__1_) );
  NOR2X1 U304 ( .A(n72), .B(n46), .Y(ab_2__19_) );
  NOR2X1 U305 ( .A(n71), .B(n46), .Y(ab_2__18_) );
  NOR2X1 U306 ( .A(n70), .B(n46), .Y(ab_2__17_) );
  NOR2X1 U307 ( .A(n69), .B(n47), .Y(ab_2__16_) );
  NOR2X1 U308 ( .A(n67), .B(n47), .Y(ab_2__15_) );
  NOR2X1 U309 ( .A(n66), .B(n47), .Y(ab_2__14_) );
  NOR2X1 U310 ( .A(n65), .B(n47), .Y(ab_2__13_) );
  NOR2X1 U311 ( .A(n64), .B(n47), .Y(ab_2__12_) );
  NOR2X1 U312 ( .A(n63), .B(n47), .Y(ab_2__11_) );
  NOR2X1 U313 ( .A(n62), .B(n47), .Y(ab_2__10_) );
  NOR2X1 U314 ( .A(n37), .B(n47), .Y(ab_2__0_) );
  NOR2X1 U315 ( .A(n46), .B(n82), .Y(ab_29__2_) );
  NOR2X1 U316 ( .A(n42), .B(n82), .Y(ab_29__1_) );
  NOR2X1 U317 ( .A(n37), .B(n82), .Y(ab_29__0_) );
  NOR2X1 U318 ( .A(n50), .B(n81), .Y(ab_28__3_) );
  NOR2X1 U319 ( .A(n46), .B(n81), .Y(ab_28__2_) );
  NOR2X1 U320 ( .A(n42), .B(n81), .Y(ab_28__1_) );
  NOR2X1 U321 ( .A(n37), .B(n81), .Y(ab_28__0_) );
  NOR2X1 U322 ( .A(n55), .B(n80), .Y(ab_27__4_) );
  NOR2X1 U323 ( .A(n50), .B(n80), .Y(ab_27__3_) );
  NOR2X1 U324 ( .A(n46), .B(n80), .Y(ab_27__2_) );
  NOR2X1 U325 ( .A(n42), .B(n80), .Y(ab_27__1_) );
  NOR2X1 U326 ( .A(n37), .B(n80), .Y(ab_27__0_) );
  NOR2X1 U327 ( .A(n56), .B(n79), .Y(ab_26__5_) );
  NOR2X1 U328 ( .A(n55), .B(n79), .Y(ab_26__4_) );
  NOR2X1 U329 ( .A(n50), .B(n79), .Y(ab_26__3_) );
  NOR2X1 U330 ( .A(n46), .B(n79), .Y(ab_26__2_) );
  NOR2X1 U331 ( .A(n42), .B(n79), .Y(ab_26__1_) );
  NOR2X1 U332 ( .A(n37), .B(n79), .Y(ab_26__0_) );
  NOR2X1 U333 ( .A(n57), .B(n78), .Y(ab_25__6_) );
  NOR2X1 U334 ( .A(n56), .B(n78), .Y(ab_25__5_) );
  NOR2X1 U335 ( .A(n55), .B(n78), .Y(ab_25__4_) );
  NOR2X1 U336 ( .A(n50), .B(n78), .Y(ab_25__3_) );
  NOR2X1 U337 ( .A(n46), .B(n78), .Y(ab_25__2_) );
  NOR2X1 U338 ( .A(n42), .B(n78), .Y(ab_25__1_) );
  NOR2X1 U339 ( .A(n37), .B(n78), .Y(ab_25__0_) );
  NOR2X1 U340 ( .A(n58), .B(n77), .Y(ab_24__7_) );
  NOR2X1 U341 ( .A(n57), .B(n77), .Y(ab_24__6_) );
  NOR2X1 U342 ( .A(n56), .B(n77), .Y(ab_24__5_) );
  NOR2X1 U343 ( .A(n55), .B(n77), .Y(ab_24__4_) );
  NOR2X1 U344 ( .A(n50), .B(n77), .Y(ab_24__3_) );
  NOR2X1 U345 ( .A(n46), .B(n77), .Y(ab_24__2_) );
  NOR2X1 U346 ( .A(n42), .B(n77), .Y(ab_24__1_) );
  NOR2X1 U347 ( .A(n37), .B(n77), .Y(ab_24__0_) );
  NOR2X1 U348 ( .A(n59), .B(n76), .Y(ab_23__8_) );
  NOR2X1 U349 ( .A(n58), .B(n76), .Y(ab_23__7_) );
  NOR2X1 U350 ( .A(n57), .B(n76), .Y(ab_23__6_) );
  NOR2X1 U351 ( .A(n56), .B(n76), .Y(ab_23__5_) );
  NOR2X1 U352 ( .A(n55), .B(n76), .Y(ab_23__4_) );
  NOR2X1 U353 ( .A(n50), .B(n76), .Y(ab_23__3_) );
  NOR2X1 U354 ( .A(n46), .B(n76), .Y(ab_23__2_) );
  NOR2X1 U355 ( .A(n42), .B(n76), .Y(ab_23__1_) );
  NOR2X1 U356 ( .A(n37), .B(n76), .Y(ab_23__0_) );
  NOR2X1 U357 ( .A(n60), .B(n75), .Y(ab_22__9_) );
  NOR2X1 U358 ( .A(n59), .B(n75), .Y(ab_22__8_) );
  NOR2X1 U359 ( .A(n58), .B(n75), .Y(ab_22__7_) );
  NOR2X1 U360 ( .A(n57), .B(n75), .Y(ab_22__6_) );
  NOR2X1 U361 ( .A(n56), .B(n75), .Y(ab_22__5_) );
  NOR2X1 U362 ( .A(n55), .B(n75), .Y(ab_22__4_) );
  NOR2X1 U363 ( .A(n50), .B(n75), .Y(ab_22__3_) );
  NOR2X1 U364 ( .A(n46), .B(n75), .Y(ab_22__2_) );
  NOR2X1 U365 ( .A(n42), .B(n75), .Y(ab_22__1_) );
  NOR2X1 U366 ( .A(n37), .B(n75), .Y(ab_22__0_) );
  NOR2X1 U367 ( .A(n60), .B(n74), .Y(ab_21__9_) );
  NOR2X1 U368 ( .A(n59), .B(n74), .Y(ab_21__8_) );
  NOR2X1 U369 ( .A(n58), .B(n74), .Y(ab_21__7_) );
  NOR2X1 U370 ( .A(n57), .B(n74), .Y(ab_21__6_) );
  NOR2X1 U371 ( .A(n56), .B(n74), .Y(ab_21__5_) );
  NOR2X1 U372 ( .A(n55), .B(n74), .Y(ab_21__4_) );
  NOR2X1 U373 ( .A(n50), .B(n74), .Y(ab_21__3_) );
  NOR2X1 U374 ( .A(n46), .B(n74), .Y(ab_21__2_) );
  NOR2X1 U375 ( .A(n42), .B(n74), .Y(ab_21__1_) );
  NOR2X1 U376 ( .A(n62), .B(n74), .Y(ab_21__10_) );
  NOR2X1 U377 ( .A(n37), .B(n74), .Y(ab_21__0_) );
  NOR2X1 U378 ( .A(n60), .B(n73), .Y(ab_20__9_) );
  NOR2X1 U379 ( .A(n59), .B(n73), .Y(ab_20__8_) );
  NOR2X1 U380 ( .A(n58), .B(n73), .Y(ab_20__7_) );
  NOR2X1 U381 ( .A(n57), .B(n73), .Y(ab_20__6_) );
  NOR2X1 U382 ( .A(n56), .B(n73), .Y(ab_20__5_) );
  NOR2X1 U383 ( .A(n55), .B(n73), .Y(ab_20__4_) );
  NOR2X1 U384 ( .A(n50), .B(n73), .Y(ab_20__3_) );
  NOR2X1 U385 ( .A(n46), .B(n73), .Y(ab_20__2_) );
  NOR2X1 U386 ( .A(n41), .B(n73), .Y(ab_20__1_) );
  NOR2X1 U387 ( .A(n63), .B(n73), .Y(ab_20__11_) );
  NOR2X1 U388 ( .A(n62), .B(n73), .Y(ab_20__10_) );
  NOR2X1 U389 ( .A(n39), .B(n73), .Y(ab_20__0_) );
  NOR2X1 U390 ( .A(n60), .B(n42), .Y(ab_1__9_) );
  NOR2X1 U391 ( .A(n59), .B(n42), .Y(ab_1__8_) );
  NOR2X1 U392 ( .A(n58), .B(n42), .Y(ab_1__7_) );
  NOR2X1 U393 ( .A(n57), .B(n42), .Y(ab_1__6_) );
  NOR2X1 U394 ( .A(n56), .B(n42), .Y(ab_1__5_) );
  NOR2X1 U395 ( .A(n54), .B(n42), .Y(ab_1__4_) );
  NOR2X1 U396 ( .A(n49), .B(n42), .Y(ab_1__3_) );
  NOR2X1 U397 ( .A(n68), .B(n42), .Y(ab_1__30_) );
  NOR2X1 U398 ( .A(n45), .B(n42), .Y(ab_1__2_) );
  NOR2X1 U399 ( .A(n82), .B(n42), .Y(ab_1__29_) );
  NOR2X1 U400 ( .A(n81), .B(n42), .Y(ab_1__28_) );
  NOR2X1 U401 ( .A(n80), .B(n42), .Y(ab_1__27_) );
  NOR2X1 U402 ( .A(n79), .B(n42), .Y(ab_1__26_) );
  NOR2X1 U403 ( .A(n78), .B(n42), .Y(ab_1__25_) );
  NOR2X1 U404 ( .A(n77), .B(n42), .Y(ab_1__24_) );
  NOR2X1 U405 ( .A(n76), .B(n42), .Y(ab_1__23_) );
  NOR2X1 U406 ( .A(n75), .B(n42), .Y(ab_1__22_) );
  NOR2X1 U407 ( .A(n74), .B(n42), .Y(ab_1__21_) );
  NOR2X1 U408 ( .A(n73), .B(n42), .Y(ab_1__20_) );
  NOR2X1 U409 ( .A(n72), .B(n42), .Y(ab_1__19_) );
  NOR2X1 U410 ( .A(n71), .B(n42), .Y(ab_1__18_) );
  NOR2X1 U411 ( .A(n70), .B(n42), .Y(ab_1__17_) );
  NOR2X1 U412 ( .A(n69), .B(n42), .Y(ab_1__16_) );
  NOR2X1 U413 ( .A(n67), .B(n43), .Y(ab_1__15_) );
  NOR2X1 U414 ( .A(n66), .B(n43), .Y(ab_1__14_) );
  NOR2X1 U415 ( .A(n65), .B(n43), .Y(ab_1__13_) );
  NOR2X1 U416 ( .A(n64), .B(n43), .Y(ab_1__12_) );
  NOR2X1 U417 ( .A(n63), .B(n43), .Y(ab_1__11_) );
  NOR2X1 U418 ( .A(n62), .B(n43), .Y(ab_1__10_) );
  NOR2X1 U419 ( .A(n38), .B(n43), .Y(ab_1__0_) );
  NOR2X1 U420 ( .A(n60), .B(n72), .Y(ab_19__9_) );
  NOR2X1 U421 ( .A(n59), .B(n72), .Y(ab_19__8_) );
  NOR2X1 U422 ( .A(n58), .B(n72), .Y(ab_19__7_) );
  NOR2X1 U423 ( .A(n57), .B(n72), .Y(ab_19__6_) );
  NOR2X1 U424 ( .A(n56), .B(n72), .Y(ab_19__5_) );
  NOR2X1 U425 ( .A(n54), .B(n72), .Y(ab_19__4_) );
  NOR2X1 U426 ( .A(n49), .B(n72), .Y(ab_19__3_) );
  NOR2X1 U427 ( .A(n45), .B(n72), .Y(ab_19__2_) );
  NOR2X1 U428 ( .A(n41), .B(n72), .Y(ab_19__1_) );
  NOR2X1 U429 ( .A(n64), .B(n72), .Y(ab_19__12_) );
  NOR2X1 U430 ( .A(n63), .B(n72), .Y(ab_19__11_) );
  NOR2X1 U431 ( .A(n62), .B(n72), .Y(ab_19__10_) );
  NOR2X1 U432 ( .A(n37), .B(n72), .Y(ab_19__0_) );
  NOR2X1 U433 ( .A(n60), .B(n71), .Y(ab_18__9_) );
  NOR2X1 U434 ( .A(n59), .B(n71), .Y(ab_18__8_) );
  NOR2X1 U435 ( .A(n58), .B(n71), .Y(ab_18__7_) );
  NOR2X1 U436 ( .A(n57), .B(n71), .Y(ab_18__6_) );
  NOR2X1 U437 ( .A(n56), .B(n71), .Y(ab_18__5_) );
  NOR2X1 U438 ( .A(n54), .B(n71), .Y(ab_18__4_) );
  NOR2X1 U439 ( .A(n49), .B(n71), .Y(ab_18__3_) );
  NOR2X1 U440 ( .A(n45), .B(n71), .Y(ab_18__2_) );
  NOR2X1 U441 ( .A(n41), .B(n71), .Y(ab_18__1_) );
  NOR2X1 U442 ( .A(n65), .B(n71), .Y(ab_18__13_) );
  NOR2X1 U443 ( .A(n64), .B(n71), .Y(ab_18__12_) );
  NOR2X1 U444 ( .A(n63), .B(n71), .Y(ab_18__11_) );
  NOR2X1 U445 ( .A(n62), .B(n71), .Y(ab_18__10_) );
  NOR2X1 U446 ( .A(n39), .B(n71), .Y(ab_18__0_) );
  NOR2X1 U447 ( .A(n60), .B(n70), .Y(ab_17__9_) );
  NOR2X1 U448 ( .A(n59), .B(n70), .Y(ab_17__8_) );
  NOR2X1 U449 ( .A(n58), .B(n70), .Y(ab_17__7_) );
  NOR2X1 U450 ( .A(n57), .B(n70), .Y(ab_17__6_) );
  NOR2X1 U451 ( .A(n56), .B(n70), .Y(ab_17__5_) );
  NOR2X1 U452 ( .A(n54), .B(n70), .Y(ab_17__4_) );
  NOR2X1 U453 ( .A(n49), .B(n70), .Y(ab_17__3_) );
  NOR2X1 U454 ( .A(n45), .B(n70), .Y(ab_17__2_) );
  NOR2X1 U455 ( .A(n41), .B(n70), .Y(ab_17__1_) );
  NOR2X1 U456 ( .A(n66), .B(n70), .Y(ab_17__14_) );
  NOR2X1 U457 ( .A(n65), .B(n70), .Y(ab_17__13_) );
  NOR2X1 U458 ( .A(n64), .B(n70), .Y(ab_17__12_) );
  NOR2X1 U459 ( .A(n63), .B(n70), .Y(ab_17__11_) );
  NOR2X1 U460 ( .A(n62), .B(n70), .Y(ab_17__10_) );
  NOR2X1 U461 ( .A(n37), .B(n70), .Y(ab_17__0_) );
  NOR2X1 U462 ( .A(n61), .B(n69), .Y(ab_16__9_) );
  NOR2X1 U463 ( .A(n59), .B(n69), .Y(ab_16__8_) );
  NOR2X1 U464 ( .A(n58), .B(n69), .Y(ab_16__7_) );
  NOR2X1 U465 ( .A(n57), .B(n69), .Y(ab_16__6_) );
  NOR2X1 U466 ( .A(n56), .B(n69), .Y(ab_16__5_) );
  NOR2X1 U467 ( .A(n54), .B(n69), .Y(ab_16__4_) );
  NOR2X1 U468 ( .A(n49), .B(n69), .Y(ab_16__3_) );
  NOR2X1 U469 ( .A(n45), .B(n69), .Y(ab_16__2_) );
  NOR2X1 U470 ( .A(n41), .B(n69), .Y(ab_16__1_) );
  NOR2X1 U471 ( .A(n67), .B(n69), .Y(ab_16__15_) );
  NOR2X1 U472 ( .A(n66), .B(n69), .Y(ab_16__14_) );
  NOR2X1 U473 ( .A(n65), .B(n69), .Y(ab_16__13_) );
  NOR2X1 U474 ( .A(n64), .B(n69), .Y(ab_16__12_) );
  NOR2X1 U475 ( .A(n63), .B(n69), .Y(ab_16__11_) );
  NOR2X1 U476 ( .A(n62), .B(n69), .Y(ab_16__10_) );
  NOR2X1 U477 ( .A(n39), .B(n69), .Y(ab_16__0_) );
  NOR2X1 U478 ( .A(n61), .B(n67), .Y(ab_15__9_) );
  NOR2X1 U479 ( .A(n59), .B(n67), .Y(ab_15__8_) );
  NOR2X1 U480 ( .A(n58), .B(n67), .Y(ab_15__7_) );
  NOR2X1 U481 ( .A(n57), .B(n67), .Y(ab_15__6_) );
  NOR2X1 U482 ( .A(n56), .B(n67), .Y(ab_15__5_) );
  NOR2X1 U483 ( .A(n54), .B(n67), .Y(ab_15__4_) );
  NOR2X1 U484 ( .A(n49), .B(n67), .Y(ab_15__3_) );
  NOR2X1 U485 ( .A(n45), .B(n67), .Y(ab_15__2_) );
  NOR2X1 U486 ( .A(n41), .B(n67), .Y(ab_15__1_) );
  NOR2X1 U487 ( .A(n69), .B(n67), .Y(ab_15__16_) );
  NOR2X1 U488 ( .A(n66), .B(n67), .Y(ab_15__14_) );
  NOR2X1 U489 ( .A(n65), .B(n67), .Y(ab_15__13_) );
  NOR2X1 U490 ( .A(n64), .B(n67), .Y(ab_15__12_) );
  NOR2X1 U491 ( .A(n63), .B(n67), .Y(ab_15__11_) );
  NOR2X1 U492 ( .A(n62), .B(n67), .Y(ab_15__10_) );
  NOR2X1 U493 ( .A(n37), .B(n67), .Y(ab_15__0_) );
  NOR2X1 U494 ( .A(n61), .B(n66), .Y(ab_14__9_) );
  NOR2X1 U495 ( .A(n59), .B(n66), .Y(ab_14__8_) );
  NOR2X1 U496 ( .A(n58), .B(n66), .Y(ab_14__7_) );
  NOR2X1 U497 ( .A(n57), .B(n66), .Y(ab_14__6_) );
  NOR2X1 U498 ( .A(n56), .B(n66), .Y(ab_14__5_) );
  NOR2X1 U499 ( .A(n54), .B(n66), .Y(ab_14__4_) );
  NOR2X1 U500 ( .A(n49), .B(n66), .Y(ab_14__3_) );
  NOR2X1 U501 ( .A(n45), .B(n66), .Y(ab_14__2_) );
  NOR2X1 U502 ( .A(n41), .B(n66), .Y(ab_14__1_) );
  NOR2X1 U503 ( .A(n70), .B(n66), .Y(ab_14__17_) );
  NOR2X1 U504 ( .A(n69), .B(n66), .Y(ab_14__16_) );
  NOR2X1 U505 ( .A(n67), .B(n66), .Y(ab_14__15_) );
  NOR2X1 U506 ( .A(n65), .B(n66), .Y(ab_14__13_) );
  NOR2X1 U507 ( .A(n64), .B(n66), .Y(ab_14__12_) );
  NOR2X1 U508 ( .A(n63), .B(n66), .Y(ab_14__11_) );
  NOR2X1 U509 ( .A(n62), .B(n66), .Y(ab_14__10_) );
  NOR2X1 U510 ( .A(n37), .B(n66), .Y(ab_14__0_) );
  NOR2X1 U511 ( .A(n61), .B(n65), .Y(ab_13__9_) );
  NOR2X1 U512 ( .A(n59), .B(n65), .Y(ab_13__8_) );
  NOR2X1 U513 ( .A(n58), .B(n65), .Y(ab_13__7_) );
  NOR2X1 U514 ( .A(n57), .B(n65), .Y(ab_13__6_) );
  NOR2X1 U515 ( .A(n56), .B(n65), .Y(ab_13__5_) );
  NOR2X1 U516 ( .A(n54), .B(n65), .Y(ab_13__4_) );
  NOR2X1 U517 ( .A(n49), .B(n65), .Y(ab_13__3_) );
  NOR2X1 U518 ( .A(n45), .B(n65), .Y(ab_13__2_) );
  NOR2X1 U519 ( .A(n41), .B(n65), .Y(ab_13__1_) );
  NOR2X1 U520 ( .A(n71), .B(n65), .Y(ab_13__18_) );
  NOR2X1 U521 ( .A(n70), .B(n65), .Y(ab_13__17_) );
  NOR2X1 U522 ( .A(n69), .B(n65), .Y(ab_13__16_) );
  NOR2X1 U523 ( .A(n67), .B(n65), .Y(ab_13__15_) );
  NOR2X1 U524 ( .A(n66), .B(n65), .Y(ab_13__14_) );
  NOR2X1 U525 ( .A(n64), .B(n65), .Y(ab_13__12_) );
  NOR2X1 U526 ( .A(n63), .B(n65), .Y(ab_13__11_) );
  NOR2X1 U527 ( .A(n62), .B(n65), .Y(ab_13__10_) );
  NOR2X1 U528 ( .A(n39), .B(n65), .Y(ab_13__0_) );
  NOR2X1 U529 ( .A(n61), .B(n64), .Y(ab_12__9_) );
  NOR2X1 U530 ( .A(n59), .B(n64), .Y(ab_12__8_) );
  NOR2X1 U531 ( .A(n58), .B(n64), .Y(ab_12__7_) );
  NOR2X1 U532 ( .A(n57), .B(n64), .Y(ab_12__6_) );
  NOR2X1 U533 ( .A(n56), .B(n64), .Y(ab_12__5_) );
  NOR2X1 U534 ( .A(n54), .B(n64), .Y(ab_12__4_) );
  NOR2X1 U535 ( .A(n49), .B(n64), .Y(ab_12__3_) );
  NOR2X1 U536 ( .A(n45), .B(n64), .Y(ab_12__2_) );
  NOR2X1 U537 ( .A(n41), .B(n64), .Y(ab_12__1_) );
  NOR2X1 U538 ( .A(n72), .B(n64), .Y(ab_12__19_) );
  NOR2X1 U539 ( .A(n71), .B(n64), .Y(ab_12__18_) );
  NOR2X1 U540 ( .A(n70), .B(n64), .Y(ab_12__17_) );
  NOR2X1 U541 ( .A(n69), .B(n64), .Y(ab_12__16_) );
  NOR2X1 U542 ( .A(n67), .B(n64), .Y(ab_12__15_) );
  NOR2X1 U543 ( .A(n66), .B(n64), .Y(ab_12__14_) );
  NOR2X1 U544 ( .A(n65), .B(n64), .Y(ab_12__13_) );
  NOR2X1 U545 ( .A(n63), .B(n64), .Y(ab_12__11_) );
  NOR2X1 U546 ( .A(n62), .B(n64), .Y(ab_12__10_) );
  NOR2X1 U547 ( .A(n37), .B(n64), .Y(ab_12__0_) );
  NOR2X1 U548 ( .A(n61), .B(n63), .Y(ab_11__9_) );
  NOR2X1 U549 ( .A(n59), .B(n63), .Y(ab_11__8_) );
  NOR2X1 U550 ( .A(n58), .B(n63), .Y(ab_11__7_) );
  NOR2X1 U551 ( .A(n57), .B(n63), .Y(ab_11__6_) );
  NOR2X1 U552 ( .A(n56), .B(n63), .Y(ab_11__5_) );
  NOR2X1 U553 ( .A(n54), .B(n63), .Y(ab_11__4_) );
  NOR2X1 U554 ( .A(n49), .B(n63), .Y(ab_11__3_) );
  NOR2X1 U555 ( .A(n45), .B(n63), .Y(ab_11__2_) );
  NOR2X1 U556 ( .A(n73), .B(n63), .Y(ab_11__20_) );
  NOR2X1 U557 ( .A(n41), .B(n63), .Y(ab_11__1_) );
  NOR2X1 U558 ( .A(n72), .B(n63), .Y(ab_11__19_) );
  NOR2X1 U559 ( .A(n71), .B(n63), .Y(ab_11__18_) );
  NOR2X1 U560 ( .A(n70), .B(n63), .Y(ab_11__17_) );
  NOR2X1 U561 ( .A(n69), .B(n63), .Y(ab_11__16_) );
  NOR2X1 U562 ( .A(n67), .B(n63), .Y(ab_11__15_) );
  NOR2X1 U563 ( .A(n66), .B(n63), .Y(ab_11__14_) );
  NOR2X1 U564 ( .A(n65), .B(n63), .Y(ab_11__13_) );
  NOR2X1 U565 ( .A(n64), .B(n63), .Y(ab_11__12_) );
  NOR2X1 U566 ( .A(n62), .B(n63), .Y(ab_11__10_) );
  NOR2X1 U567 ( .A(n39), .B(n63), .Y(ab_11__0_) );
  NOR2X1 U568 ( .A(n61), .B(n62), .Y(ab_10__9_) );
  NOR2X1 U569 ( .A(n59), .B(n62), .Y(ab_10__8_) );
  NOR2X1 U570 ( .A(n58), .B(n62), .Y(ab_10__7_) );
  NOR2X1 U571 ( .A(n57), .B(n62), .Y(ab_10__6_) );
  NOR2X1 U572 ( .A(n56), .B(n62), .Y(ab_10__5_) );
  NOR2X1 U573 ( .A(n54), .B(n62), .Y(ab_10__4_) );
  NOR2X1 U574 ( .A(n49), .B(n62), .Y(ab_10__3_) );
  NOR2X1 U575 ( .A(n45), .B(n62), .Y(ab_10__2_) );
  NOR2X1 U576 ( .A(n74), .B(n62), .Y(ab_10__21_) );
  NOR2X1 U577 ( .A(n73), .B(n62), .Y(ab_10__20_) );
  NOR2X1 U578 ( .A(n41), .B(n62), .Y(ab_10__1_) );
  NOR2X1 U579 ( .A(n72), .B(n62), .Y(ab_10__19_) );
  NOR2X1 U580 ( .A(n71), .B(n62), .Y(ab_10__18_) );
  NOR2X1 U581 ( .A(n70), .B(n62), .Y(ab_10__17_) );
  NOR2X1 U582 ( .A(n69), .B(n62), .Y(ab_10__16_) );
  NOR2X1 U583 ( .A(n67), .B(n62), .Y(ab_10__15_) );
  NOR2X1 U584 ( .A(n66), .B(n62), .Y(ab_10__14_) );
  NOR2X1 U585 ( .A(n65), .B(n62), .Y(ab_10__13_) );
  NOR2X1 U586 ( .A(n64), .B(n62), .Y(ab_10__12_) );
  NOR2X1 U587 ( .A(n63), .B(n62), .Y(ab_10__11_) );
  NOR2X1 U588 ( .A(n39), .B(n62), .Y(ab_10__0_) );
  NOR2X1 U589 ( .A(n61), .B(n39), .Y(ab_0__9_) );
  NOR2X1 U590 ( .A(n59), .B(n39), .Y(ab_0__8_) );
  NOR2X1 U591 ( .A(n58), .B(n39), .Y(ab_0__7_) );
  NOR2X1 U592 ( .A(n57), .B(n39), .Y(ab_0__6_) );
  NOR2X1 U593 ( .A(n56), .B(n39), .Y(ab_0__5_) );
  NOR2X1 U594 ( .A(n54), .B(n39), .Y(ab_0__4_) );
  NOR2X1 U595 ( .A(n49), .B(n39), .Y(ab_0__3_) );
  NOR2X1 U596 ( .A(n68), .B(n39), .Y(ab_0__30_) );
  NOR2X1 U597 ( .A(n45), .B(n39), .Y(ab_0__2_) );
  NOR2X1 U598 ( .A(n82), .B(n38), .Y(ab_0__29_) );
  NOR2X1 U599 ( .A(n81), .B(n38), .Y(ab_0__28_) );
  NOR2X1 U600 ( .A(n80), .B(n38), .Y(ab_0__27_) );
  NOR2X1 U601 ( .A(n79), .B(n38), .Y(ab_0__26_) );
  NOR2X1 U602 ( .A(n78), .B(n38), .Y(ab_0__25_) );
  NOR2X1 U603 ( .A(n77), .B(n38), .Y(ab_0__24_) );
  NOR2X1 U604 ( .A(n76), .B(n38), .Y(ab_0__23_) );
  NOR2X1 U605 ( .A(n75), .B(n38), .Y(ab_0__22_) );
  NOR2X1 U606 ( .A(n74), .B(n38), .Y(ab_0__21_) );
  NOR2X1 U607 ( .A(n73), .B(n38), .Y(ab_0__20_) );
  NOR2X1 U608 ( .A(n41), .B(n38), .Y(ab_0__1_) );
  NOR2X1 U609 ( .A(n72), .B(n38), .Y(ab_0__19_) );
  NOR2X1 U610 ( .A(n71), .B(n38), .Y(ab_0__18_) );
  NOR2X1 U611 ( .A(n70), .B(n38), .Y(ab_0__17_) );
  NOR2X1 U612 ( .A(n69), .B(n39), .Y(ab_0__16_) );
  NOR2X1 U613 ( .A(n67), .B(n37), .Y(ab_0__15_) );
  NOR2X1 U614 ( .A(n66), .B(n39), .Y(ab_0__14_) );
  NOR2X1 U615 ( .A(n65), .B(n39), .Y(ab_0__13_) );
  NOR2X1 U616 ( .A(n64), .B(n37), .Y(ab_0__12_) );
  NOR2X1 U617 ( .A(n63), .B(n39), .Y(ab_0__11_) );
  NOR2X1 U618 ( .A(n62), .B(n39), .Y(ab_0__10_) );
endmodule


module square_root_finder ( rst, clk, in, sqrt );
  input [15:0] in;
  output [31:0] sqrt;
  input rst, clk;
  wire   n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, cat_0_, N30, N31, N32, N33, N34, N35, N36, N37, N38,
         N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N83, N84,
         N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98,
         N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, N292, n118, n120,
         n121, n122, n123, n124, n125, n126, n127, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n1490, n1510, n1520, n1530, n1540,
         n1550, n1560, n1570, n1580, n1590, n1600, n1610, n1620, n1630, n1640,
         n1650, n1660, n1670, n1680, n1690, n1700, n1710, n1720, n1730, n1740,
         n1750, n1760, n1770, n1780, n1790, n180, n181, n182, n184, n185,
         n1860, n1870, n1880, n1890, n1900, n1910, n1920, n1930, n1940, n1950,
         n1960, n1970, n1980, n1990, n2000, n2010, n2020, n2030, n2040, n2050,
         n2060, n2070, n2080, n2090, n2100, n2110, n2120, n2130, n2140, n2150,
         n2160, n2170, n2180, n2190, n2200, n2210, n2220, n2230, n2240, n2250,
         n2260, n2270, n2280, n2290, n2300, n2310, n2320, n2330, n2340, n2350,
         n2360, n2370, n2380, n2390, n2400, n2410, n2420, n2430, n2440, n2460,
         n2470, n248, n249, n250, n251, n252, n253, n254, n255, n258, n261,
         n264, n267, n270, n273, n276, n279, n282, n285, n288, n291, n294,
         n297, n300, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         N1480, N1470, N1460, N1450, N1440, N1430, N1420, N1410, N1400, N1390,
         N1380, N1370, N1360, N1350, N1340, N1330, N1320, N1310, N1300, N1290,
         N128, N1270, N1260, N1250, N1240, N1230, N1220, N1210, N1200, N119,
         N1180, N117, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72,
         N71, N70, N69, N68, N67, N66, N65, N64, N63, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n366, n367, n369, n371, n373, n375, n377, n378, n379, n381, n382,
         n383, n384, n386, n388, n390, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475;
  wire   [1:0] state;
  wire   [31:0] up;
  wire   [31:0] low;
  wire   [31:13] sub_51_carry;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111;

  square_root_finder_DW01_add_0 add_80 ( .A({1'b0, sqrt[30:0]}), .B({1'b0, 
        low[30:0]}), .CI(1'b0), .SUM({N247, N246, N245, N244, N243, N242, N241, 
        N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, 
        SYNOPSYS_UNCONNECTED__0}), .CO() );
  square_root_finder_DW01_add_1 add_73 ( .A({1'b0, up[30:0]}), .B({1'b0, 
        sqrt[30:0]}), .CI(1'b0), .SUM({N216, N215, N214, N213, N212, N211, 
        N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, 
        N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        N186, SYNOPSYS_UNCONNECTED__1}), .CO() );
  square_root_finder_DW02_mult_2 mult_31 ( .A({1'b0, sqrt[30:0]}), .B({1'b0, 
        sqrt[30:0]}), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45}) );
  square_root_finder_DW02_mult_1 mult_33 ( .A({1'b0, sqrt[30:0]}), .B({1'b0, 
        sqrt[30:0]}), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, 
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, N1480, N1470, N1460, N1450, N1440, N1430, 
        N1420, N1410, N1400, N1390, N1380, N1370, N1360, N1350, N1340, N1330, 
        N1320, N1310, N1300, N1290, N128, N1270, N1260, N1250, N1240, N1230, 
        N1220, N1210, N1200, N119, N1180, N117}) );
  square_root_finder_DW01_sub_1 sub_33 ( .A({1'b0, 1'b0, 1'b0, 1'b0, in, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({N1480, N1470, N1460, N1450, N1440, N1430, N1420, N1410, N1400, 
        N1390, N1380, N1370, N1360, N1350, N1340, N1330, N1320, N1310, N1300, 
        N1290, N128, N1270, N1260, N1250, N1240, N1230, N1220, N1210, N1200, 
        N119, N1180, N117}), .CI(1'b0), .DIFF({N179, N178, N177, N176, N175, 
        N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, SYNOPSYS_UNCONNECTED__78}), .CO() );
  square_root_finder_DW02_mult_0 mult_51 ( .A({1'b0, sqrt[30:0]}), .B({1'b0, 
        sqrt[30:0]}), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, N82, N81, N80, N79, N78, N77, N76, N75, N74, 
        N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N93, N92, N91, 
        N90, N89, N88, N87, N86, N85, N84, N83, SYNOPSYS_UNCONNECTED__111}) );
  DFFRHQX1 up_reg_30_ ( .D(n2460), .CK(clk), .RN(rst), .Q(up[30]) );
  DFFRHQX1 up_reg_28_ ( .D(n248), .CK(clk), .RN(rst), .Q(up[28]) );
  DFFRHQX1 up_reg_29_ ( .D(n2470), .CK(clk), .RN(rst), .Q(up[29]) );
  DFFRHQX1 low_reg_30_ ( .D(n184), .CK(clk), .RN(rst), .Q(low[30]) );
  DFFRHQX1 low_reg_28_ ( .D(n1860), .CK(clk), .RN(rst), .Q(low[28]) );
  DFFRHQX1 low_reg_29_ ( .D(n185), .CK(clk), .RN(rst), .Q(low[29]) );
  DFFRHQX1 up_reg_24_ ( .D(n252), .CK(clk), .RN(rst), .Q(up[24]) );
  DFFRHQX1 up_reg_25_ ( .D(n251), .CK(clk), .RN(rst), .Q(up[25]) );
  DFFRHQX1 up_reg_26_ ( .D(n250), .CK(clk), .RN(rst), .Q(up[26]) );
  DFFRHQX1 up_reg_27_ ( .D(n249), .CK(clk), .RN(rst), .Q(up[27]) );
  DFFRHQX1 low_reg_24_ ( .D(n1900), .CK(clk), .RN(rst), .Q(low[24]) );
  DFFRHQX1 low_reg_25_ ( .D(n1890), .CK(clk), .RN(rst), .Q(low[25]) );
  DFFRHQX1 low_reg_26_ ( .D(n1880), .CK(clk), .RN(rst), .Q(low[26]) );
  DFFRHQX1 low_reg_27_ ( .D(n1870), .CK(clk), .RN(rst), .Q(low[27]) );
  DFFRHQX1 cat_reg_0_ ( .D(n310), .CK(clk), .RN(rst), .Q(cat_0_) );
  DFFRHQX1 state_reg_0_ ( .D(n311), .CK(clk), .RN(rst), .Q(state[0]) );
  DFFRHQX1 up_reg_22_ ( .D(n254), .CK(clk), .RN(rst), .Q(up[22]) );
  DFFRHQX1 up_reg_23_ ( .D(n253), .CK(clk), .RN(rst), .Q(up[23]) );
  DFFRHQX1 low_reg_19_ ( .D(n1950), .CK(clk), .RN(rst), .Q(low[19]) );
  DFFRHQX1 low_reg_20_ ( .D(n1940), .CK(clk), .RN(rst), .Q(low[20]) );
  DFFRHQX1 low_reg_21_ ( .D(n1930), .CK(clk), .RN(rst), .Q(low[21]) );
  DFFRHQX1 low_reg_22_ ( .D(n1920), .CK(clk), .RN(rst), .Q(low[22]) );
  DFFRHQX1 low_reg_23_ ( .D(n1910), .CK(clk), .RN(rst), .Q(low[23]) );
  DFFSRHQX1 up_reg_20_ ( .D(n258), .CK(clk), .SN(n319), .RN(n335), .Q(up[20])
         );
  DFFRHQX1 low_reg_15_ ( .D(n1990), .CK(clk), .RN(rst), .Q(low[15]) );
  DFFRHQX1 low_reg_16_ ( .D(n1980), .CK(clk), .RN(rst), .Q(low[16]) );
  DFFRHQX1 low_reg_17_ ( .D(n1970), .CK(clk), .RN(rst), .Q(low[17]) );
  DFFRHQX1 low_reg_18_ ( .D(n1960), .CK(clk), .RN(rst), .Q(low[18]) );
  DFFSRHQX1 up_reg_16_ ( .D(n270), .CK(clk), .SN(n323), .RN(n339), .Q(up[16])
         );
  DFFSRHQX1 up_reg_17_ ( .D(n267), .CK(clk), .SN(n322), .RN(n338), .Q(up[17])
         );
  DFFSRHQX1 up_reg_18_ ( .D(n264), .CK(clk), .SN(n321), .RN(n337), .Q(up[18])
         );
  DFFSRHQX1 up_reg_19_ ( .D(n261), .CK(clk), .SN(n320), .RN(n336), .Q(up[19])
         );
  DFFRHQX1 low_reg_11_ ( .D(n2030), .CK(clk), .RN(rst), .Q(low[11]) );
  DFFRHQX1 low_reg_12_ ( .D(n2020), .CK(clk), .RN(rst), .Q(low[12]) );
  DFFRHQX1 low_reg_13_ ( .D(n2010), .CK(clk), .RN(rst), .Q(low[13]) );
  DFFRHQX1 low_reg_14_ ( .D(n2000), .CK(clk), .RN(rst), .Q(low[14]) );
  DFFSRHQX1 up_reg_12_ ( .D(n282), .CK(clk), .SN(n327), .RN(n343), .Q(up[12])
         );
  DFFSRHQX1 up_reg_13_ ( .D(n279), .CK(clk), .SN(n326), .RN(n342), .Q(up[13])
         );
  DFFSRHQX1 up_reg_14_ ( .D(n276), .CK(clk), .SN(n325), .RN(n341), .Q(up[14])
         );
  DFFSRHQX1 up_reg_15_ ( .D(n273), .CK(clk), .SN(n324), .RN(n340), .Q(up[15])
         );
  DFFRHQX1 low_reg_7_ ( .D(n2070), .CK(clk), .RN(rst), .Q(low[7]) );
  DFFRHQX1 low_reg_8_ ( .D(n2060), .CK(clk), .RN(rst), .Q(low[8]) );
  DFFRHQX1 low_reg_9_ ( .D(n2050), .CK(clk), .RN(rst), .Q(low[9]) );
  DFFRHQX1 low_reg_10_ ( .D(n2040), .CK(clk), .RN(rst), .Q(low[10]) );
  DFFSRHQX1 up_reg_7_ ( .D(n297), .CK(clk), .SN(n332), .RN(n348), .Q(up[7]) );
  DFFSRHQX1 up_reg_8_ ( .D(n294), .CK(clk), .SN(n331), .RN(n347), .Q(up[8]) );
  DFFSRHQX1 up_reg_9_ ( .D(n291), .CK(clk), .SN(n330), .RN(n346), .Q(up[9]) );
  DFFSRHQX1 up_reg_10_ ( .D(n288), .CK(clk), .SN(n329), .RN(n345), .Q(up[10])
         );
  DFFSRHQX1 up_reg_11_ ( .D(n285), .CK(clk), .SN(n328), .RN(n344), .Q(up[11])
         );
  DFFRHQX1 up_reg_3_ ( .D(n305), .CK(clk), .RN(rst), .Q(up[3]) );
  DFFRHQX1 up_reg_4_ ( .D(n304), .CK(clk), .RN(rst), .Q(up[4]) );
  DFFRHQX1 up_reg_5_ ( .D(n303), .CK(clk), .RN(rst), .Q(up[5]) );
  DFFRHQX1 low_reg_2_ ( .D(n2120), .CK(clk), .RN(rst), .Q(low[2]) );
  DFFRHQX1 low_reg_3_ ( .D(n2110), .CK(clk), .RN(rst), .Q(low[3]) );
  DFFRHQX1 low_reg_4_ ( .D(n2100), .CK(clk), .RN(rst), .Q(low[4]) );
  DFFRHQX1 low_reg_5_ ( .D(n2090), .CK(clk), .RN(rst), .Q(low[5]) );
  DFFRHQX1 low_reg_6_ ( .D(n2080), .CK(clk), .RN(rst), .Q(low[6]) );
  DFFSRHQX1 up_reg_6_ ( .D(n300), .CK(clk), .SN(n333), .RN(n349), .Q(up[6]) );
  DFFRHQX1 low_reg_0_ ( .D(n2140), .CK(clk), .RN(rst), .Q(low[0]) );
  DFFRHQX1 up_reg_0_ ( .D(n308), .CK(clk), .RN(rst), .Q(up[0]) );
  DFFRHQX1 up_reg_1_ ( .D(n307), .CK(clk), .RN(rst), .Q(up[1]) );
  DFFRHQX1 up_reg_2_ ( .D(n306), .CK(clk), .RN(rst), .Q(up[2]) );
  DFFRHQX1 low_reg_1_ ( .D(n2130), .CK(clk), .RN(rst), .Q(low[1]) );
  DFFRHQX1 g_reg_30_ ( .D(n2150), .CK(clk), .RN(rst), .Q(n482) );
  DFFRHQX1 g_reg_24_ ( .D(n2210), .CK(clk), .RN(rst), .Q(n488) );
  DFFRHQX1 g_reg_25_ ( .D(n2200), .CK(clk), .RN(rst), .Q(n487) );
  DFFRHQX1 g_reg_26_ ( .D(n2190), .CK(clk), .RN(rst), .Q(n486) );
  DFFRHQX1 g_reg_27_ ( .D(n2180), .CK(clk), .RN(rst), .Q(n485) );
  DFFRHQX1 g_reg_28_ ( .D(n2170), .CK(clk), .RN(rst), .Q(n484) );
  DFFRHQX1 g_reg_29_ ( .D(n2160), .CK(clk), .RN(rst), .Q(n483) );
  DFFRHQX1 g_reg_13_ ( .D(n2320), .CK(clk), .RN(rst), .Q(n498) );
  DFFRHQX1 g_reg_14_ ( .D(n2310), .CK(clk), .RN(rst), .Q(n497) );
  DFFRHQX1 g_reg_15_ ( .D(n2300), .CK(clk), .RN(rst), .Q(sqrt[15]) );
  DFFRHQX1 g_reg_16_ ( .D(n2290), .CK(clk), .RN(rst), .Q(n496) );
  DFFRHQX1 g_reg_17_ ( .D(n2280), .CK(clk), .RN(rst), .Q(n495) );
  DFFRHQX1 g_reg_18_ ( .D(n2270), .CK(clk), .RN(rst), .Q(n494) );
  DFFRHQX1 g_reg_19_ ( .D(n2260), .CK(clk), .RN(rst), .Q(n493) );
  DFFRHQX1 g_reg_20_ ( .D(n2250), .CK(clk), .RN(rst), .Q(n492) );
  DFFRHQX1 g_reg_21_ ( .D(n2240), .CK(clk), .RN(rst), .Q(n491) );
  DFFRHQX1 g_reg_22_ ( .D(n2230), .CK(clk), .RN(rst), .Q(n490) );
  DFFRHQX1 g_reg_23_ ( .D(n2220), .CK(clk), .RN(rst), .Q(n489) );
  DFFRHQX1 g_reg_6_ ( .D(n2390), .CK(clk), .RN(rst), .Q(sqrt[6]) );
  DFFRHQX1 g_reg_7_ ( .D(n2380), .CK(clk), .RN(rst), .Q(n501) );
  DFFRHQX1 g_reg_8_ ( .D(n2370), .CK(clk), .RN(rst), .Q(sqrt[8]) );
  DFFRHQX1 g_reg_9_ ( .D(n2360), .CK(clk), .RN(rst), .Q(sqrt[9]) );
  DFFRHQX1 g_reg_10_ ( .D(n2350), .CK(clk), .RN(rst), .Q(sqrt[10]) );
  DFFRHQX1 g_reg_11_ ( .D(n2340), .CK(clk), .RN(rst), .Q(n500) );
  DFFRHQX1 g_reg_12_ ( .D(n2330), .CK(clk), .RN(rst), .Q(n499) );
  DFFRHQX1 g_reg_0_ ( .D(n309), .CK(clk), .RN(rst), .Q(n506) );
  DFFRHQX1 g_reg_1_ ( .D(n2440), .CK(clk), .RN(rst), .Q(n505) );
  DFFRHQX1 g_reg_2_ ( .D(n2430), .CK(clk), .RN(rst), .Q(n504) );
  DFFRHQX1 g_reg_3_ ( .D(n2420), .CK(clk), .RN(rst), .Q(n503) );
  DFFRHQX1 g_reg_4_ ( .D(n2410), .CK(clk), .RN(rst), .Q(n502) );
  DFFRHQX1 g_reg_5_ ( .D(n2400), .CK(clk), .RN(rst), .Q(sqrt[5]) );
  DFFSRXL up_reg_21_ ( .D(n255), .CK(clk), .SN(n318), .RN(n334), .Q(up[21]), 
        .QN(n467) );
  DFFRXL state_reg_1_ ( .D(state[0]), .CK(clk), .RN(rst), .Q(state[1]), .QN(
        n443) );
  INVX1 U306 ( .A(1'b1), .Y(sqrt[31]) );
  NAND2X1 U308 ( .A(n442), .B(n126), .Y(n314) );
  NAND2X1 U309 ( .A(N292), .B(n1510), .Y(n315) );
  NAND2X1 U310 ( .A(N292), .B(n182), .Y(n316) );
  NOR4X1 U311 ( .A(N155), .B(N154), .C(N153), .D(N152), .Y(n138) );
  NOR4X1 U312 ( .A(N91), .B(N90), .C(N89), .D(N88), .Y(n146) );
  INVX1 U313 ( .A(n1510), .Y(n367) );
  NOR2X1 U314 ( .A(n139), .B(n140), .Y(n124) );
  NAND4X1 U315 ( .A(n145), .B(n146), .C(n147), .D(n148), .Y(n139) );
  NAND4X1 U316 ( .A(n141), .B(n142), .C(n143), .D(n144), .Y(n140) );
  NOR4X1 U317 ( .A(N87), .B(N86), .C(N85), .D(N84), .Y(n145) );
  INVX1 U318 ( .A(n316), .Y(n442) );
  INVX1 U319 ( .A(n182), .Y(n366) );
  NOR4X1 U320 ( .A(N83), .B(N50), .C(N113), .D(N112), .Y(n144) );
  NAND2X1 U321 ( .A(N50), .B(n317), .Y(n123) );
  NOR4X1 U322 ( .A(N179), .B(N178), .C(N177), .D(N176), .Y(n137) );
  OAI22X1 U323 ( .A0(n121), .A1(n444), .B0(n122), .B1(n123), .Y(n310) );
  AOI211X1 U324 ( .A0(n124), .A1(n317), .B0(n125), .C0(n126), .Y(n121) );
  NAND2X1 U325 ( .A(n127), .B(n123), .Y(n125) );
  NAND4BXL U326 ( .AN(n124), .B(n350), .C(n127), .D(n129), .Y(n311) );
  AOI21X1 U327 ( .A0(n122), .A1(n440), .B0(n126), .Y(n129) );
  INVX1 U328 ( .A(n123), .Y(n440) );
  AND4X2 U329 ( .A(n130), .B(n131), .C(n132), .D(n133), .Y(n122) );
  NOR4BX1 U330 ( .AN(n138), .B(N151), .C(N149), .D(N150), .Y(n132) );
  NOR4X1 U331 ( .A(N159), .B(N158), .C(N157), .D(N156), .Y(n130) );
  NOR4X1 U332 ( .A(N163), .B(N162), .C(N161), .D(N160), .Y(n131) );
  INVX1 U333 ( .A(n381), .Y(sqrt[7]) );
  INVX1 U334 ( .A(n386), .Y(sqrt[11]) );
  INVX1 U335 ( .A(n388), .Y(sqrt[12]) );
  INVX1 U336 ( .A(n369), .Y(sqrt[0]) );
  AND4X2 U337 ( .A(n134), .B(n135), .C(n136), .D(n137), .Y(n133) );
  NOR4X1 U338 ( .A(N167), .B(N166), .C(N165), .D(N164), .Y(n134) );
  NOR4X1 U339 ( .A(N171), .B(N170), .C(N169), .D(N168), .Y(n135) );
  NOR4X1 U340 ( .A(N175), .B(N174), .C(N173), .D(N172), .Y(n136) );
  INVX1 U341 ( .A(n371), .Y(sqrt[1]) );
  INVX1 U342 ( .A(n373), .Y(sqrt[2]) );
  INVX1 U343 ( .A(n375), .Y(sqrt[3]) );
  INVX1 U344 ( .A(n377), .Y(sqrt[4]) );
  NOR4X1 U345 ( .A(N111), .B(N110), .C(N109), .D(N108), .Y(n143) );
  INVX1 U346 ( .A(n390), .Y(sqrt[13]) );
  INVX1 U347 ( .A(n392), .Y(sqrt[14]) );
  NOR4X1 U348 ( .A(N107), .B(N106), .C(N105), .D(N104), .Y(n142) );
  NOR4X1 U349 ( .A(N103), .B(N102), .C(N101), .D(N100), .Y(n141) );
  NOR4X1 U350 ( .A(N99), .B(N98), .C(N97), .D(N96), .Y(n148) );
  NOR4X1 U351 ( .A(N95), .B(N94), .C(N93), .D(N92), .Y(n147) );
  OAI21XL U352 ( .A0(N292), .A1(n475), .B0(n1530), .Y(n2160) );
  AOI22X1 U353 ( .A0(N246), .A1(n367), .B0(N215), .B1(n366), .Y(n1530) );
  OAI21XL U354 ( .A0(N292), .A1(n474), .B0(n1540), .Y(n2170) );
  AOI22X1 U355 ( .A0(N245), .A1(n367), .B0(N214), .B1(n366), .Y(n1540) );
  OAI21XL U356 ( .A0(N292), .A1(n473), .B0(n1550), .Y(n2180) );
  AOI22X1 U357 ( .A0(N244), .A1(n367), .B0(N213), .B1(n366), .Y(n1550) );
  OAI21XL U358 ( .A0(N292), .A1(n472), .B0(n1560), .Y(n2190) );
  AOI22X1 U359 ( .A0(N243), .A1(n367), .B0(N212), .B1(n366), .Y(n1560) );
  OAI21XL U360 ( .A0(N292), .A1(n471), .B0(n1570), .Y(n2200) );
  AOI22X1 U361 ( .A0(N242), .A1(n367), .B0(N211), .B1(n366), .Y(n1570) );
  OAI21XL U362 ( .A0(N292), .A1(n470), .B0(n1580), .Y(n2210) );
  AOI22X1 U363 ( .A0(N241), .A1(n367), .B0(N210), .B1(n366), .Y(n1580) );
  OAI21XL U364 ( .A0(N292), .A1(n469), .B0(n1590), .Y(n2220) );
  AOI22X1 U365 ( .A0(N240), .A1(n367), .B0(N209), .B1(n366), .Y(n1590) );
  OAI21XL U366 ( .A0(N292), .A1(n468), .B0(n1600), .Y(n2230) );
  AOI22X1 U367 ( .A0(N239), .A1(n367), .B0(N208), .B1(n366), .Y(n1600) );
  OAI21XL U368 ( .A0(N292), .A1(n466), .B0(n1610), .Y(n2240) );
  AOI22X1 U369 ( .A0(N238), .A1(n367), .B0(N207), .B1(n366), .Y(n1610) );
  OAI21XL U370 ( .A0(N292), .A1(n464), .B0(n1620), .Y(n2250) );
  AOI22X1 U371 ( .A0(N237), .A1(n367), .B0(N206), .B1(n366), .Y(n1620) );
  OAI21XL U372 ( .A0(N292), .A1(n462), .B0(n1630), .Y(n2260) );
  AOI22X1 U373 ( .A0(N236), .A1(n367), .B0(N205), .B1(n366), .Y(n1630) );
  OAI21XL U374 ( .A0(N292), .A1(n460), .B0(n1640), .Y(n2270) );
  AOI22X1 U375 ( .A0(N235), .A1(n367), .B0(N204), .B1(n366), .Y(n1640) );
  OAI21XL U376 ( .A0(N292), .A1(n458), .B0(n1650), .Y(n2280) );
  AOI22X1 U377 ( .A0(N234), .A1(n367), .B0(N203), .B1(n366), .Y(n1650) );
  OAI21XL U378 ( .A0(N292), .A1(n456), .B0(n1660), .Y(n2290) );
  AOI22X1 U379 ( .A0(N233), .A1(n367), .B0(N202), .B1(n366), .Y(n1660) );
  OAI21XL U380 ( .A0(N292), .A1(n393), .B0(n1670), .Y(n2300) );
  AOI22X1 U381 ( .A0(N232), .A1(n367), .B0(N201), .B1(n366), .Y(n1670) );
  OAI21XL U382 ( .A0(N292), .A1(n392), .B0(n1680), .Y(n2310) );
  AOI22X1 U383 ( .A0(N231), .A1(n367), .B0(N200), .B1(n366), .Y(n1680) );
  OAI21XL U384 ( .A0(N292), .A1(n390), .B0(n1690), .Y(n2320) );
  AOI22X1 U385 ( .A0(N230), .A1(n367), .B0(N199), .B1(n366), .Y(n1690) );
  OAI21XL U386 ( .A0(N292), .A1(n378), .B0(n1770), .Y(n2400) );
  AOI22X1 U387 ( .A0(N222), .A1(n367), .B0(N191), .B1(n366), .Y(n1770) );
  NAND2X1 U388 ( .A(n126), .B(n444), .Y(n1510) );
  OAI21XL U389 ( .A0(N292), .A1(n377), .B0(n1780), .Y(n2410) );
  AOI22X1 U390 ( .A0(N221), .A1(n367), .B0(N190), .B1(n366), .Y(n1780) );
  OAI21XL U391 ( .A0(N292), .A1(n375), .B0(n1790), .Y(n2420) );
  AOI22X1 U392 ( .A0(N220), .A1(n367), .B0(N189), .B1(n366), .Y(n1790) );
  OAI21XL U393 ( .A0(N292), .A1(n373), .B0(n180), .Y(n2430) );
  AOI22X1 U394 ( .A0(N219), .A1(n367), .B0(N188), .B1(n366), .Y(n180) );
  OAI21XL U395 ( .A0(N292), .A1(n371), .B0(n181), .Y(n2440) );
  AOI22X1 U396 ( .A0(N218), .A1(n367), .B0(N187), .B1(n366), .Y(n181) );
  NOR2BX1 U397 ( .AN(n127), .B(n317), .Y(N292) );
  NAND2BX1 U398 ( .AN(n315), .B(n126), .Y(n1490) );
  OAI21XL U399 ( .A0(N292), .A1(n369), .B0(n120), .Y(n309) );
  AOI22X1 U400 ( .A0(N217), .A1(n367), .B0(N186), .B1(n366), .Y(n120) );
  INVX1 U401 ( .A(sqrt[16]), .Y(n456) );
  INVX1 U402 ( .A(sqrt[17]), .Y(n458) );
  INVX1 U403 ( .A(sqrt[18]), .Y(n460) );
  INVX1 U404 ( .A(sqrt[19]), .Y(n462) );
  INVX1 U405 ( .A(sqrt[20]), .Y(n464) );
  INVX1 U406 ( .A(sqrt[21]), .Y(n466) );
  INVX1 U407 ( .A(sqrt[22]), .Y(n468) );
  INVX1 U408 ( .A(sqrt[23]), .Y(n469) );
  INVX1 U409 ( .A(sqrt[24]), .Y(n470) );
  INVX1 U410 ( .A(sqrt[25]), .Y(n471) );
  INVX1 U411 ( .A(sqrt[26]), .Y(n472) );
  INVX1 U412 ( .A(sqrt[27]), .Y(n473) );
  INVX1 U413 ( .A(sqrt[28]), .Y(n474) );
  INVX1 U414 ( .A(sqrt[29]), .Y(n475) );
  INVX1 U415 ( .A(sqrt[30]), .Y(n445) );
  ADDFX2 U416 ( .A(N78), .B(n402), .CI(sub_51_carry[27]), .CO(sub_51_carry[28]), .S(N109) );
  INVX1 U417 ( .A(in[15]), .Y(n402) );
  ADDFX2 U418 ( .A(N76), .B(n401), .CI(sub_51_carry[25]), .CO(sub_51_carry[26]), .S(N107) );
  INVX1 U419 ( .A(in[13]), .Y(n401) );
  ADDFX2 U420 ( .A(N77), .B(n425), .CI(sub_51_carry[26]), .CO(sub_51_carry[27]), .S(N108) );
  INVX1 U421 ( .A(n499), .Y(n388) );
  INVX1 U422 ( .A(n500), .Y(n386) );
  INVX1 U423 ( .A(sqrt[10]), .Y(n384) );
  INVX1 U424 ( .A(sqrt[9]), .Y(n383) );
  INVX1 U425 ( .A(sqrt[8]), .Y(n382) );
  INVX1 U426 ( .A(n501), .Y(n381) );
  INVX1 U427 ( .A(sqrt[6]), .Y(n379) );
  INVX1 U428 ( .A(sqrt[5]), .Y(n378) );
  INVX1 U429 ( .A(n502), .Y(n377) );
  INVX1 U430 ( .A(n503), .Y(n375) );
  INVX1 U431 ( .A(n504), .Y(n373) );
  INVX1 U432 ( .A(n505), .Y(n371) );
  INVX1 U433 ( .A(n506), .Y(n369) );
  INVX1 U434 ( .A(N42), .Y(n436) );
  INVX1 U435 ( .A(N43), .Y(n437) );
  BUFX3 U436 ( .A(n496), .Y(sqrt[16]) );
  BUFX3 U437 ( .A(n495), .Y(sqrt[17]) );
  BUFX3 U438 ( .A(n494), .Y(sqrt[18]) );
  BUFX3 U439 ( .A(n493), .Y(sqrt[19]) );
  BUFX3 U440 ( .A(n492), .Y(sqrt[20]) );
  BUFX3 U441 ( .A(n491), .Y(sqrt[21]) );
  BUFX3 U442 ( .A(n490), .Y(sqrt[22]) );
  BUFX3 U443 ( .A(n489), .Y(sqrt[23]) );
  ADDFX2 U444 ( .A(N67), .B(n420), .CI(sub_51_carry[16]), .CO(sub_51_carry[17]), .S(N98) );
  ADDFX2 U445 ( .A(N68), .B(n397), .CI(sub_51_carry[17]), .CO(sub_51_carry[18]), .S(N99) );
  INVX1 U446 ( .A(in[5]), .Y(n397) );
  ADDFX2 U447 ( .A(N69), .B(n421), .CI(sub_51_carry[18]), .CO(sub_51_carry[19]), .S(N100) );
  ADDFX2 U448 ( .A(N70), .B(n398), .CI(sub_51_carry[19]), .CO(sub_51_carry[20]), .S(N101) );
  INVX1 U449 ( .A(in[7]), .Y(n398) );
  ADDFX2 U450 ( .A(N71), .B(n422), .CI(sub_51_carry[20]), .CO(sub_51_carry[21]), .S(N102) );
  ADDFX2 U451 ( .A(N72), .B(n399), .CI(sub_51_carry[21]), .CO(sub_51_carry[22]), .S(N103) );
  INVX1 U452 ( .A(in[9]), .Y(n399) );
  ADDFX2 U453 ( .A(N73), .B(n423), .CI(sub_51_carry[22]), .CO(sub_51_carry[23]), .S(N104) );
  ADDFX2 U454 ( .A(N74), .B(n400), .CI(sub_51_carry[23]), .CO(sub_51_carry[24]), .S(N105) );
  INVX1 U455 ( .A(in[11]), .Y(n400) );
  ADDFX2 U456 ( .A(N75), .B(n424), .CI(sub_51_carry[24]), .CO(sub_51_carry[25]), .S(N106) );
  INVX1 U457 ( .A(sqrt[15]), .Y(n393) );
  INVX1 U458 ( .A(n497), .Y(n392) );
  INVX1 U459 ( .A(n498), .Y(n390) );
  INVX1 U460 ( .A(N44), .Y(n438) );
  INVX1 U461 ( .A(N45), .Y(n439) );
  INVX1 U462 ( .A(N36), .Y(n430) );
  INVX1 U463 ( .A(N37), .Y(n431) );
  INVX1 U464 ( .A(N38), .Y(n432) );
  INVX1 U465 ( .A(N39), .Y(n433) );
  INVX1 U466 ( .A(N40), .Y(n434) );
  INVX1 U467 ( .A(N41), .Y(n435) );
  BUFX3 U468 ( .A(n488), .Y(sqrt[24]) );
  BUFX3 U469 ( .A(n487), .Y(sqrt[25]) );
  BUFX3 U470 ( .A(n486), .Y(sqrt[26]) );
  BUFX3 U471 ( .A(n485), .Y(sqrt[27]) );
  BUFX3 U472 ( .A(n484), .Y(sqrt[28]) );
  ADDFX2 U473 ( .A(N64), .B(n441), .CI(sub_51_carry[13]), .CO(sub_51_carry[14]), .S(N95) );
  ADDFX2 U474 ( .A(N65), .B(n395), .CI(sub_51_carry[14]), .CO(sub_51_carry[15]), .S(N96) );
  INVX1 U475 ( .A(in[2]), .Y(n395) );
  ADDFX2 U476 ( .A(N66), .B(n396), .CI(sub_51_carry[15]), .CO(sub_51_carry[16]), .S(N97) );
  INVX1 U477 ( .A(in[3]), .Y(n396) );
  BUFX3 U478 ( .A(n483), .Y(sqrt[29]) );
  BUFX3 U479 ( .A(n482), .Y(sqrt[30]) );
  INVX1 U480 ( .A(N32), .Y(n426) );
  INVX1 U481 ( .A(N33), .Y(n427) );
  INVX1 U482 ( .A(N34), .Y(n428) );
  INVX1 U483 ( .A(N35), .Y(n429) );
  OAI21XL U484 ( .A0(N292), .A1(n445), .B0(n1520), .Y(n2150) );
  AOI22X1 U485 ( .A0(N247), .A1(n367), .B0(N216), .B1(n366), .Y(n1520) );
  OAI21XL U486 ( .A0(N292), .A1(n388), .B0(n1700), .Y(n2330) );
  AOI22X1 U487 ( .A0(N229), .A1(n367), .B0(N198), .B1(n366), .Y(n1700) );
  OAI21XL U488 ( .A0(N292), .A1(n386), .B0(n1710), .Y(n2340) );
  AOI22X1 U489 ( .A0(N228), .A1(n367), .B0(N197), .B1(n366), .Y(n1710) );
  OAI21XL U490 ( .A0(N292), .A1(n384), .B0(n1720), .Y(n2350) );
  AOI22X1 U491 ( .A0(N227), .A1(n367), .B0(N196), .B1(n366), .Y(n1720) );
  OAI21XL U492 ( .A0(N292), .A1(n383), .B0(n1730), .Y(n2360) );
  AOI22X1 U493 ( .A0(N226), .A1(n367), .B0(N195), .B1(n366), .Y(n1730) );
  OAI21XL U494 ( .A0(N292), .A1(n382), .B0(n1740), .Y(n2370) );
  AOI22X1 U495 ( .A0(N225), .A1(n367), .B0(N194), .B1(n366), .Y(n1740) );
  OAI21XL U496 ( .A0(N292), .A1(n381), .B0(n1750), .Y(n2380) );
  AOI22X1 U497 ( .A0(N224), .A1(n367), .B0(N193), .B1(n366), .Y(n1750) );
  OAI21XL U498 ( .A0(N292), .A1(n379), .B0(n1760), .Y(n2390) );
  AOI22X1 U499 ( .A0(N223), .A1(n367), .B0(N192), .B1(n366), .Y(n1760) );
  OAI222XL U500 ( .A0(n314), .A1(n466), .B0(n350), .B1(n402), .C0(n442), .C1(
        n467), .Y(n255) );
  OAI222XL U501 ( .A0(n314), .A1(n464), .B0(n350), .B1(n425), .C0(n442), .C1(
        n465), .Y(n258) );
  INVX1 U502 ( .A(up[20]), .Y(n465) );
  OAI222XL U503 ( .A0(n314), .A1(n462), .B0(n350), .B1(n401), .C0(n442), .C1(
        n463), .Y(n261) );
  INVX1 U504 ( .A(up[19]), .Y(n463) );
  OAI222XL U505 ( .A0(n314), .A1(n460), .B0(n350), .B1(n424), .C0(n442), .C1(
        n461), .Y(n264) );
  INVX1 U506 ( .A(up[18]), .Y(n461) );
  OAI222XL U507 ( .A0(n314), .A1(n458), .B0(n350), .B1(n400), .C0(n442), .C1(
        n459), .Y(n267) );
  INVX1 U508 ( .A(up[17]), .Y(n459) );
  OAI222XL U509 ( .A0(n314), .A1(n456), .B0(n350), .B1(n423), .C0(n442), .C1(
        n457), .Y(n270) );
  INVX1 U510 ( .A(up[16]), .Y(n457) );
  OAI222XL U511 ( .A0(n314), .A1(n393), .B0(n350), .B1(n399), .C0(n442), .C1(
        n455), .Y(n273) );
  INVX1 U512 ( .A(up[15]), .Y(n455) );
  OAI222XL U513 ( .A0(n314), .A1(n392), .B0(n350), .B1(n422), .C0(n442), .C1(
        n454), .Y(n276) );
  INVX1 U514 ( .A(up[14]), .Y(n454) );
  OAI222XL U515 ( .A0(n314), .A1(n390), .B0(n398), .B1(n350), .C0(n442), .C1(
        n453), .Y(n279) );
  INVX1 U516 ( .A(up[13]), .Y(n453) );
  OAI222XL U517 ( .A0(n314), .A1(n388), .B0(n350), .B1(n421), .C0(n442), .C1(
        n452), .Y(n282) );
  INVX1 U518 ( .A(up[12]), .Y(n452) );
  OAI222XL U519 ( .A0(n314), .A1(n386), .B0(n350), .B1(n397), .C0(n442), .C1(
        n451), .Y(n285) );
  INVX1 U520 ( .A(up[11]), .Y(n451) );
  OAI222XL U521 ( .A0(n314), .A1(n384), .B0(n350), .B1(n420), .C0(n442), .C1(
        n450), .Y(n288) );
  INVX1 U522 ( .A(up[10]), .Y(n450) );
  OAI222XL U523 ( .A0(n314), .A1(n383), .B0(n350), .B1(n396), .C0(n442), .C1(
        n449), .Y(n291) );
  INVX1 U524 ( .A(up[9]), .Y(n449) );
  OAI222XL U525 ( .A0(n314), .A1(n382), .B0(n350), .B1(n395), .C0(n442), .C1(
        n448), .Y(n294) );
  INVX1 U526 ( .A(up[8]), .Y(n448) );
  OAI222XL U527 ( .A0(n314), .A1(n381), .B0(n350), .B1(n441), .C0(n442), .C1(
        n447), .Y(n297) );
  INVX1 U528 ( .A(up[7]), .Y(n447) );
  OAI222XL U529 ( .A0(n314), .A1(n379), .B0(n350), .B1(n394), .C0(n442), .C1(
        n446), .Y(n300) );
  INVX1 U530 ( .A(up[6]), .Y(n446) );
  NOR2X1 U531 ( .A(n443), .B(state[0]), .Y(n126) );
  NAND2X1 U532 ( .A(state[1]), .B(state[0]), .Y(n127) );
  NAND2X1 U533 ( .A(cat_0_), .B(n126), .Y(n182) );
  OAI2BB2X1 U534 ( .B0(n314), .B1(n475), .A0N(up[29]), .A1N(n316), .Y(n2470)
         );
  OAI2BB2X1 U535 ( .B0(n1490), .B1(n475), .A0N(low[29]), .A1N(n315), .Y(n185)
         );
  OAI2BB2X1 U536 ( .B0(n314), .B1(n474), .A0N(up[28]), .A1N(n316), .Y(n248) );
  OAI2BB2X1 U537 ( .B0(n1490), .B1(n474), .A0N(low[28]), .A1N(n315), .Y(n1860)
         );
  OAI2BB2X1 U538 ( .B0(n314), .B1(n473), .A0N(up[27]), .A1N(n316), .Y(n249) );
  OAI2BB2X1 U539 ( .B0(n1490), .B1(n473), .A0N(low[27]), .A1N(n315), .Y(n1870)
         );
  OAI2BB2X1 U540 ( .B0(n314), .B1(n472), .A0N(up[26]), .A1N(n316), .Y(n250) );
  OAI2BB2X1 U541 ( .B0(n1490), .B1(n472), .A0N(low[26]), .A1N(n315), .Y(n1880)
         );
  OAI2BB2X1 U542 ( .B0(n314), .B1(n471), .A0N(up[25]), .A1N(n316), .Y(n251) );
  OAI2BB2X1 U543 ( .B0(n1490), .B1(n471), .A0N(low[25]), .A1N(n315), .Y(n1890)
         );
  OAI2BB2X1 U544 ( .B0(n314), .B1(n470), .A0N(up[24]), .A1N(n316), .Y(n252) );
  OAI2BB2X1 U545 ( .B0(n1490), .B1(n470), .A0N(low[24]), .A1N(n315), .Y(n1900)
         );
  OAI2BB2X1 U546 ( .B0(n314), .B1(n469), .A0N(up[23]), .A1N(n316), .Y(n253) );
  OAI2BB2X1 U547 ( .B0(n1490), .B1(n469), .A0N(low[23]), .A1N(n315), .Y(n1910)
         );
  OAI2BB2X1 U548 ( .B0(n314), .B1(n468), .A0N(up[22]), .A1N(n316), .Y(n254) );
  OAI2BB2X1 U549 ( .B0(n1490), .B1(n468), .A0N(low[22]), .A1N(n315), .Y(n1920)
         );
  OAI2BB2X1 U550 ( .B0(n1490), .B1(n466), .A0N(low[21]), .A1N(n315), .Y(n1930)
         );
  OAI2BB2X1 U551 ( .B0(n1490), .B1(n464), .A0N(low[20]), .A1N(n315), .Y(n1940)
         );
  OAI2BB2X1 U552 ( .B0(n1490), .B1(n462), .A0N(low[19]), .A1N(n315), .Y(n1950)
         );
  OAI2BB2X1 U553 ( .B0(n1490), .B1(n460), .A0N(low[18]), .A1N(n315), .Y(n1960)
         );
  OAI2BB2X1 U554 ( .B0(n1490), .B1(n458), .A0N(low[17]), .A1N(n315), .Y(n1970)
         );
  OAI2BB2X1 U555 ( .B0(n1490), .B1(n456), .A0N(low[16]), .A1N(n315), .Y(n1980)
         );
  OAI2BB2X1 U556 ( .B0(n388), .B1(n1490), .A0N(low[12]), .A1N(n315), .Y(n2020)
         );
  OAI2BB2X1 U557 ( .B0(n386), .B1(n1490), .A0N(low[11]), .A1N(n315), .Y(n2030)
         );
  OAI2BB2X1 U558 ( .B0(n384), .B1(n1490), .A0N(low[10]), .A1N(n315), .Y(n2040)
         );
  OAI2BB2X1 U559 ( .B0(n383), .B1(n1490), .A0N(low[9]), .A1N(n315), .Y(n2050)
         );
  OAI2BB2X1 U560 ( .B0(n382), .B1(n1490), .A0N(low[8]), .A1N(n315), .Y(n2060)
         );
  OAI2BB2X1 U561 ( .B0(n381), .B1(n1490), .A0N(low[7]), .A1N(n315), .Y(n2070)
         );
  OAI2BB2X1 U562 ( .B0(n379), .B1(n1490), .A0N(low[6]), .A1N(n315), .Y(n2080)
         );
  OAI2BB2X1 U563 ( .B0(n378), .B1(n1490), .A0N(low[5]), .A1N(n315), .Y(n2090)
         );
  OAI2BB2X1 U564 ( .B0(n1490), .B1(n393), .A0N(low[15]), .A1N(n315), .Y(n1990)
         );
  OAI2BB2X1 U565 ( .B0(n1490), .B1(n392), .A0N(low[14]), .A1N(n315), .Y(n2000)
         );
  OAI2BB2X1 U566 ( .B0(n1490), .B1(n390), .A0N(low[13]), .A1N(n315), .Y(n2010)
         );
  OAI2BB2X1 U567 ( .B0(n314), .B1(n378), .A0N(up[5]), .A1N(n316), .Y(n303) );
  OAI2BB2X1 U568 ( .B0(n377), .B1(n1490), .A0N(low[4]), .A1N(n315), .Y(n2100)
         );
  OAI2BB2X1 U569 ( .B0(n314), .B1(n377), .A0N(up[4]), .A1N(n316), .Y(n304) );
  OAI2BB2X1 U570 ( .B0(n375), .B1(n1490), .A0N(low[3]), .A1N(n315), .Y(n2110)
         );
  OAI2BB2X1 U571 ( .B0(n314), .B1(n375), .A0N(up[3]), .A1N(n316), .Y(n305) );
  OAI2BB2X1 U572 ( .B0(n373), .B1(n1490), .A0N(low[2]), .A1N(n315), .Y(n2120)
         );
  OAI2BB2X1 U573 ( .B0(n314), .B1(n373), .A0N(up[2]), .A1N(n316), .Y(n306) );
  OAI2BB2X1 U574 ( .B0(n371), .B1(n1490), .A0N(low[1]), .A1N(n315), .Y(n2130)
         );
  OAI2BB2X1 U575 ( .B0(n314), .B1(n371), .A0N(up[1]), .A1N(n316), .Y(n307) );
  OAI2BB2X1 U576 ( .B0(n314), .B1(n445), .A0N(up[30]), .A1N(n316), .Y(n2460)
         );
  OAI2BB2X1 U577 ( .B0(n1490), .B1(n445), .A0N(low[30]), .A1N(n315), .Y(n184)
         );
  OAI2BB2X1 U578 ( .B0(n369), .B1(n1490), .A0N(low[0]), .A1N(n315), .Y(n2140)
         );
  OAI2BB2X1 U579 ( .B0(n314), .B1(n369), .A0N(up[0]), .A1N(n316), .Y(n308) );
  INVX1 U580 ( .A(cat_0_), .Y(n444) );
  AND2X2 U581 ( .A(state[0]), .B(n443), .Y(n317) );
  BUFX3 U582 ( .A(n118), .Y(n350) );
  NAND2BX1 U583 ( .AN(state[0]), .B(n443), .Y(n118) );
  OR2X2 U584 ( .A(rst), .B(n402), .Y(n318) );
  OR2X2 U585 ( .A(rst), .B(n425), .Y(n319) );
  OR2X2 U586 ( .A(rst), .B(n401), .Y(n320) );
  OR2X2 U587 ( .A(rst), .B(n424), .Y(n321) );
  OR2X2 U588 ( .A(rst), .B(n400), .Y(n322) );
  OR2X2 U589 ( .A(rst), .B(n423), .Y(n323) );
  OR2X2 U590 ( .A(rst), .B(n399), .Y(n324) );
  OR2X2 U591 ( .A(rst), .B(n422), .Y(n325) );
  OR2X2 U592 ( .A(rst), .B(n398), .Y(n326) );
  OR2X2 U593 ( .A(rst), .B(n421), .Y(n327) );
  OR2X2 U594 ( .A(rst), .B(n397), .Y(n328) );
  OR2X2 U595 ( .A(rst), .B(n420), .Y(n329) );
  OR2X2 U596 ( .A(rst), .B(n396), .Y(n330) );
  OR2X2 U597 ( .A(rst), .B(n395), .Y(n331) );
  OR2X2 U598 ( .A(rst), .B(n441), .Y(n332) );
  OR2X2 U599 ( .A(rst), .B(n394), .Y(n333) );
  OR2X2 U600 ( .A(rst), .B(in[15]), .Y(n334) );
  OR2X2 U601 ( .A(rst), .B(in[14]), .Y(n335) );
  OR2X2 U602 ( .A(rst), .B(in[13]), .Y(n336) );
  OR2X2 U603 ( .A(rst), .B(in[12]), .Y(n337) );
  OR2X2 U604 ( .A(rst), .B(in[11]), .Y(n338) );
  OR2X2 U605 ( .A(rst), .B(in[10]), .Y(n339) );
  OR2X2 U606 ( .A(rst), .B(in[9]), .Y(n340) );
  OR2X2 U607 ( .A(rst), .B(in[8]), .Y(n341) );
  OR2X2 U608 ( .A(rst), .B(in[7]), .Y(n342) );
  OR2X2 U609 ( .A(rst), .B(in[6]), .Y(n343) );
  OR2X2 U610 ( .A(rst), .B(in[5]), .Y(n344) );
  OR2X2 U611 ( .A(rst), .B(in[4]), .Y(n345) );
  OR2X2 U612 ( .A(rst), .B(in[3]), .Y(n346) );
  OR2X2 U613 ( .A(rst), .B(in[2]), .Y(n347) );
  OR2X2 U614 ( .A(rst), .B(in[1]), .Y(n348) );
  OR2X2 U615 ( .A(rst), .B(in[0]), .Y(n349) );
  INVX1 U616 ( .A(in[1]), .Y(n441) );
  INVX1 U617 ( .A(in[0]), .Y(n394) );
  INVX1 U618 ( .A(in[4]), .Y(n420) );
  INVX1 U619 ( .A(in[6]), .Y(n421) );
  INVX1 U620 ( .A(in[8]), .Y(n422) );
  INVX1 U621 ( .A(in[10]), .Y(n423) );
  INVX1 U622 ( .A(in[12]), .Y(n424) );
  INVX1 U623 ( .A(in[14]), .Y(n425) );
  XNOR2X1 U626 ( .A(N82), .B(sub_51_carry[31]), .Y(N113) );
  OR2X1 U627 ( .A(N81), .B(sub_51_carry[30]), .Y(sub_51_carry[31]) );
  XNOR2X1 U628 ( .A(sub_51_carry[30]), .B(N81), .Y(N112) );
  OR2X1 U629 ( .A(N80), .B(sub_51_carry[29]), .Y(sub_51_carry[30]) );
  XNOR2X1 U630 ( .A(sub_51_carry[29]), .B(N80), .Y(N111) );
  OR2X1 U631 ( .A(N79), .B(sub_51_carry[28]), .Y(sub_51_carry[29]) );
  XNOR2X1 U632 ( .A(sub_51_carry[28]), .B(N79), .Y(N110) );
  OR2X1 U633 ( .A(n394), .B(N63), .Y(sub_51_carry[13]) );
  XNOR2X1 U634 ( .A(N63), .B(n394), .Y(N94) );
  NAND2BX1 U635 ( .AN(N30), .B(in[0]), .Y(n404) );
  AOI2BB1X1 U636 ( .A0N(n404), .A1N(N31), .B0(in[1]), .Y(n403) );
  AOI221X1 U637 ( .A0(N32), .A1(n395), .B0(N31), .B1(n404), .C0(n403), .Y(n405) );
  AOI221X1 U638 ( .A0(in[3]), .A1(n427), .B0(in[2]), .B1(n426), .C0(n405), .Y(
        n406) );
  AOI221X1 U639 ( .A0(N34), .A1(n420), .B0(N33), .B1(n396), .C0(n406), .Y(n407) );
  AOI221X1 U640 ( .A0(in[5]), .A1(n429), .B0(in[4]), .B1(n428), .C0(n407), .Y(
        n408) );
  AOI221X1 U641 ( .A0(N36), .A1(n421), .B0(N35), .B1(n397), .C0(n408), .Y(n409) );
  AOI221X1 U642 ( .A0(in[7]), .A1(n431), .B0(in[6]), .B1(n430), .C0(n409), .Y(
        n410) );
  AOI221X1 U643 ( .A0(N38), .A1(n422), .B0(N37), .B1(n398), .C0(n410), .Y(n411) );
  AOI221X1 U644 ( .A0(in[9]), .A1(n433), .B0(in[8]), .B1(n432), .C0(n411), .Y(
        n412) );
  AOI221X1 U645 ( .A0(N40), .A1(n423), .B0(N39), .B1(n399), .C0(n412), .Y(n413) );
  AOI221X1 U646 ( .A0(in[11]), .A1(n435), .B0(in[10]), .B1(n434), .C0(n413), 
        .Y(n414) );
  AOI221X1 U647 ( .A0(N42), .A1(n424), .B0(N41), .B1(n400), .C0(n414), .Y(n415) );
  AOI221X1 U648 ( .A0(in[13]), .A1(n437), .B0(in[12]), .B1(n436), .C0(n415), 
        .Y(n416) );
  AOI221X1 U649 ( .A0(N44), .A1(n425), .B0(N43), .B1(n401), .C0(n416), .Y(n417) );
  AOI221X1 U650 ( .A0(in[15]), .A1(n439), .B0(in[14]), .B1(n438), .C0(n417), 
        .Y(n418) );
  AOI211X1 U651 ( .A0(N45), .A1(n402), .B0(N46), .C0(n418), .Y(n419) );
  NOR4BX1 U652 ( .AN(n419), .B(N49), .C(N47), .D(N48), .Y(N50) );
endmodule

