
module square_root_finder ( rst, clk, in, sqrt );
  input [15:0] in;
  output [31:0] sqrt;
  input rst, clk;
  wire   N34, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, n42, n74, n75, n76, n77, n820,
         n830, n840, n850, n890, n900, n910, n920, n940, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n1440, n1450, n1460, n1470, n1480, n1490, n1500, n1510;
  wire   [28:14] sub_45_carry;

  DFFHQX1 inx_reg_27_ ( .D(in[15]), .CK(rst), .Q(N94) );
  DFFHQX1 inx_reg_23_ ( .D(in[11]), .CK(rst), .Q(N90) );
  DFFHQX1 inx_reg_19_ ( .D(in[7]), .CK(rst), .Q(N86) );
  DFFHQX1 inx_reg_15_ ( .D(in[3]), .CK(rst), .Q(N82) );
  DFFHQX1 inx_reg_25_ ( .D(in[13]), .CK(rst), .Q(N92) );
  DFFHQX1 inx_reg_21_ ( .D(in[9]), .CK(rst), .Q(N88) );
  DFFHQX1 inx_reg_17_ ( .D(in[5]), .CK(rst), .Q(N84) );
  DFFHQX1 inx_reg_26_ ( .D(in[14]), .CK(rst), .Q(N93) );
  DFFHQX1 inx_reg_22_ ( .D(in[10]), .CK(rst), .Q(N89) );
  DFFHQX1 inx_reg_18_ ( .D(in[6]), .CK(rst), .Q(N85) );
  DFFHQX1 inx_reg_14_ ( .D(in[2]), .CK(rst), .Q(N81) );
  DFFHQX1 inx_reg_24_ ( .D(in[12]), .CK(rst), .Q(N91) );
  DFFHQX1 inx_reg_20_ ( .D(in[8]), .CK(rst), .Q(N87) );
  DFFHQX1 inx_reg_16_ ( .D(in[4]), .CK(rst), .Q(N83) );
  DFFHQX1 inx_reg_13_ ( .D(in[1]), .CK(rst), .Q(N80) );
  DFFHQX1 inx_reg_12_ ( .D(in[0]), .CK(rst), .Q(N79) );
  DFFHQX1 sqrt_reg_31_ ( .D(n132), .CK(clk), .Q(sqrt[31]) );
  DFFHQX1 sqrt_reg_30_ ( .D(n131), .CK(clk), .Q(sqrt[30]) );
  DFFHQX1 sqrt_reg_29_ ( .D(n130), .CK(clk), .Q(sqrt[29]) );
  DFFHQX1 sqrt_reg_28_ ( .D(n129), .CK(clk), .Q(sqrt[28]) );
  DFFHQX1 sqrt_reg_27_ ( .D(n128), .CK(clk), .Q(sqrt[27]) );
  DFFHQX1 sqrt_reg_26_ ( .D(n127), .CK(clk), .Q(sqrt[26]) );
  DFFHQX1 sqrt_reg_25_ ( .D(n126), .CK(clk), .Q(sqrt[25]) );
  DFFHQX1 sqrt_reg_24_ ( .D(n125), .CK(clk), .Q(sqrt[24]) );
  DFFHQX1 sqrt_reg_23_ ( .D(n124), .CK(clk), .Q(sqrt[23]) );
  DFFHQX1 sqrt_reg_22_ ( .D(n123), .CK(clk), .Q(sqrt[22]) );
  DFFHQX1 sqrt_reg_21_ ( .D(n122), .CK(clk), .Q(sqrt[21]) );
  DFFHQX1 sqrt_reg_20_ ( .D(n121), .CK(clk), .Q(sqrt[20]) );
  DFFHQX1 sqrt_reg_19_ ( .D(n120), .CK(clk), .Q(sqrt[19]) );
  DFFHQX1 sqrt_reg_18_ ( .D(n119), .CK(clk), .Q(sqrt[18]) );
  DFFHQX1 sqrt_reg_17_ ( .D(n118), .CK(clk), .Q(sqrt[17]) );
  DFFHQX1 sqrt_reg_16_ ( .D(n117), .CK(clk), .Q(sqrt[16]) );
  DFFHQX1 sqrt_reg_15_ ( .D(n116), .CK(clk), .Q(sqrt[15]) );
  DFFHQX1 sqrt_reg_14_ ( .D(n115), .CK(clk), .Q(sqrt[14]) );
  DFFHQX1 sqrt_reg_13_ ( .D(n114), .CK(clk), .Q(sqrt[13]) );
  DFFHQX1 sqrt_reg_12_ ( .D(n113), .CK(clk), .Q(sqrt[12]) );
  DFFHQX1 sqrt_reg_11_ ( .D(n112), .CK(clk), .Q(sqrt[11]) );
  DFFHQX1 sqrt_reg_10_ ( .D(n111), .CK(clk), .Q(sqrt[10]) );
  DFFHQX1 sqrt_reg_9_ ( .D(n110), .CK(clk), .Q(sqrt[9]) );
  DFFHQX1 sqrt_reg_8_ ( .D(n109), .CK(clk), .Q(sqrt[8]) );
  DFFHQX1 sqrt_reg_7_ ( .D(n108), .CK(clk), .Q(sqrt[7]) );
  DFFHQX1 sqrt_reg_6_ ( .D(n107), .CK(clk), .Q(sqrt[6]) );
  DFFHQX1 sqrt_reg_5_ ( .D(n106), .CK(clk), .Q(sqrt[5]) );
  DFFHQX1 sqrt_reg_4_ ( .D(n105), .CK(clk), .Q(sqrt[4]) );
  DFFHQX1 sqrt_reg_3_ ( .D(n104), .CK(clk), .Q(sqrt[3]) );
  DFFHQX1 sqrt_reg_2_ ( .D(n103), .CK(clk), .Q(sqrt[2]) );
  DFFHQX1 sqrt_reg_1_ ( .D(n102), .CK(clk), .Q(sqrt[1]) );
  DFFHQX1 sqrt_reg_0_ ( .D(n101), .CK(clk), .Q(sqrt[0]) );
  OR3XL U138 ( .A(n99), .B(N90), .C(N89), .Y(n940) );
  OR3XL U139 ( .A(n100), .B(N82), .C(N81), .Y(n95) );
  OR3XL U140 ( .A(n98), .B(N86), .C(N85), .Y(n96) );
  OR3XL U141 ( .A(n940), .B(N92), .C(N91), .Y(n97) );
  OR3XL U142 ( .A(n95), .B(N84), .C(N83), .Y(n98) );
  OR3XL U143 ( .A(n96), .B(N88), .C(N87), .Y(n99) );
  OR2X2 U144 ( .A(N80), .B(N79), .Y(n100) );
  INVX1 U145 ( .A(n42), .Y(n134) );
  NOR4BX1 U146 ( .AN(sub_45_carry[28]), .B(N158), .C(N157), .D(N156), .Y(n840)
         );
  NAND4X1 U147 ( .A(n820), .B(n830), .C(n840), .D(n850), .Y(n76) );
  AND2X2 U148 ( .A(sub_45_carry[28]), .B(n1510), .Y(n850) );
  NOR4X1 U149 ( .A(N151), .B(N150), .C(N149), .D(N148), .Y(n820) );
  NOR4X1 U150 ( .A(N155), .B(N154), .C(N153), .D(N152), .Y(n830) );
  INVX1 U151 ( .A(n1510), .Y(N34) );
  OAI22X1 U152 ( .A0(n74), .A1(n75), .B0(n76), .B1(n77), .Y(n42) );
  NAND2X1 U153 ( .A(N34), .B(n890), .Y(n75) );
  AND2X2 U154 ( .A(sqrt[0]), .B(n134), .Y(n101) );
  AND2X2 U155 ( .A(sqrt[1]), .B(n134), .Y(n102) );
  AND2X2 U156 ( .A(sqrt[2]), .B(n134), .Y(n103) );
  AND2X2 U157 ( .A(sqrt[3]), .B(n134), .Y(n104) );
  AND2X2 U158 ( .A(sqrt[4]), .B(n134), .Y(n105) );
  AND2X2 U159 ( .A(sqrt[5]), .B(n134), .Y(n106) );
  AND2X2 U160 ( .A(sqrt[6]), .B(n134), .Y(n107) );
  AND2X2 U161 ( .A(sqrt[7]), .B(n134), .Y(n108) );
  AND2X2 U162 ( .A(sqrt[8]), .B(n134), .Y(n109) );
  AND2X2 U163 ( .A(sqrt[9]), .B(n134), .Y(n110) );
  AND2X2 U164 ( .A(sqrt[10]), .B(n134), .Y(n111) );
  AND2X2 U165 ( .A(sqrt[11]), .B(n134), .Y(n112) );
  AND2X2 U166 ( .A(sqrt[12]), .B(n134), .Y(n113) );
  AND2X2 U167 ( .A(sqrt[13]), .B(n134), .Y(n114) );
  AND2X2 U168 ( .A(sqrt[14]), .B(n134), .Y(n115) );
  AND2X2 U169 ( .A(sqrt[15]), .B(n134), .Y(n116) );
  AND2X2 U170 ( .A(sqrt[16]), .B(n134), .Y(n117) );
  AND2X2 U171 ( .A(sqrt[17]), .B(n134), .Y(n118) );
  AND2X2 U172 ( .A(sqrt[18]), .B(n134), .Y(n119) );
  AND2X2 U173 ( .A(sqrt[19]), .B(n134), .Y(n120) );
  AND2X2 U174 ( .A(sqrt[20]), .B(n134), .Y(n121) );
  AND2X2 U175 ( .A(sqrt[21]), .B(n134), .Y(n122) );
  AND2X2 U176 ( .A(sqrt[22]), .B(n134), .Y(n123) );
  AND2X2 U177 ( .A(sqrt[23]), .B(n134), .Y(n124) );
  AND2X2 U178 ( .A(sqrt[24]), .B(n134), .Y(n125) );
  AND2X2 U179 ( .A(sqrt[25]), .B(n134), .Y(n126) );
  AND2X2 U180 ( .A(sqrt[26]), .B(n134), .Y(n127) );
  AND2X2 U181 ( .A(sqrt[27]), .B(n134), .Y(n128) );
  AND2X2 U182 ( .A(sqrt[28]), .B(n134), .Y(n129) );
  AND2X2 U183 ( .A(sqrt[29]), .B(n134), .Y(n130) );
  AND2X2 U184 ( .A(sqrt[30]), .B(n134), .Y(n131) );
  AND2X2 U185 ( .A(sqrt[31]), .B(n134), .Y(n132) );
  NOR3X1 U186 ( .A(n97), .B(N94), .C(N93), .Y(n1510) );
  NOR4X1 U187 ( .A(N82), .B(N81), .C(N80), .D(N79), .Y(n890) );
  NAND3X1 U188 ( .A(n910), .B(n920), .C(n900), .Y(n74) );
  NOR4X1 U189 ( .A(N94), .B(N93), .C(N92), .D(N91), .Y(n920) );
  NOR4X1 U190 ( .A(N86), .B(N85), .C(N84), .D(N83), .Y(n900) );
  NOR4X1 U191 ( .A(N90), .B(N89), .C(N88), .D(N87), .Y(n910) );
  OR2X2 U192 ( .A(N79), .B(n133), .Y(n77) );
  OR4X2 U193 ( .A(N147), .B(N146), .C(N145), .D(N144), .Y(n133) );
  INVX1 U194 ( .A(N79), .Y(n135) );
  INVX1 U195 ( .A(N80), .Y(n136) );
  INVX1 U196 ( .A(N87), .Y(n143) );
  INVX1 U197 ( .A(N91), .Y(n1470) );
  INVX1 U198 ( .A(N83), .Y(n139) );
  INVX1 U199 ( .A(N85), .Y(n141) );
  INVX1 U200 ( .A(N89), .Y(n1450) );
  INVX1 U201 ( .A(N81), .Y(n137) );
  INVX1 U202 ( .A(N93), .Y(n1490) );
  INVX1 U203 ( .A(N84), .Y(n140) );
  INVX1 U204 ( .A(N88), .Y(n1440) );
  INVX1 U205 ( .A(N92), .Y(n1480) );
  INVX1 U206 ( .A(N86), .Y(n142) );
  INVX1 U207 ( .A(N90), .Y(n1460) );
  INVX1 U208 ( .A(N82), .Y(n138) );
  INVX1 U209 ( .A(N94), .Y(n1500) );
  AND2X1 U210 ( .A(sub_45_carry[27]), .B(n1500), .Y(sub_45_carry[28]) );
  XOR2X1 U211 ( .A(n1500), .B(sub_45_carry[27]), .Y(N158) );
  AND2X1 U212 ( .A(sub_45_carry[26]), .B(n1490), .Y(sub_45_carry[27]) );
  XOR2X1 U213 ( .A(n1490), .B(sub_45_carry[26]), .Y(N157) );
  AND2X1 U214 ( .A(sub_45_carry[25]), .B(n1480), .Y(sub_45_carry[26]) );
  XOR2X1 U215 ( .A(n1480), .B(sub_45_carry[25]), .Y(N156) );
  AND2X1 U216 ( .A(sub_45_carry[24]), .B(n1470), .Y(sub_45_carry[25]) );
  XOR2X1 U217 ( .A(n1470), .B(sub_45_carry[24]), .Y(N155) );
  AND2X1 U218 ( .A(sub_45_carry[23]), .B(n1460), .Y(sub_45_carry[24]) );
  XOR2X1 U219 ( .A(n1460), .B(sub_45_carry[23]), .Y(N154) );
  AND2X1 U220 ( .A(sub_45_carry[22]), .B(n1450), .Y(sub_45_carry[23]) );
  XOR2X1 U221 ( .A(n1450), .B(sub_45_carry[22]), .Y(N153) );
  AND2X1 U222 ( .A(sub_45_carry[21]), .B(n1440), .Y(sub_45_carry[22]) );
  XOR2X1 U223 ( .A(n1440), .B(sub_45_carry[21]), .Y(N152) );
  AND2X1 U224 ( .A(sub_45_carry[20]), .B(n143), .Y(sub_45_carry[21]) );
  XOR2X1 U225 ( .A(n143), .B(sub_45_carry[20]), .Y(N151) );
  AND2X1 U226 ( .A(sub_45_carry[19]), .B(n142), .Y(sub_45_carry[20]) );
  XOR2X1 U227 ( .A(n142), .B(sub_45_carry[19]), .Y(N150) );
  AND2X1 U228 ( .A(sub_45_carry[18]), .B(n141), .Y(sub_45_carry[19]) );
  XOR2X1 U229 ( .A(n141), .B(sub_45_carry[18]), .Y(N149) );
  AND2X1 U230 ( .A(sub_45_carry[17]), .B(n140), .Y(sub_45_carry[18]) );
  XOR2X1 U231 ( .A(n140), .B(sub_45_carry[17]), .Y(N148) );
  AND2X1 U232 ( .A(sub_45_carry[16]), .B(n139), .Y(sub_45_carry[17]) );
  XOR2X1 U233 ( .A(n139), .B(sub_45_carry[16]), .Y(N147) );
  AND2X1 U234 ( .A(sub_45_carry[15]), .B(n138), .Y(sub_45_carry[16]) );
  XOR2X1 U235 ( .A(n138), .B(sub_45_carry[15]), .Y(N146) );
  AND2X1 U236 ( .A(sub_45_carry[14]), .B(n137), .Y(sub_45_carry[15]) );
  XOR2X1 U237 ( .A(n137), .B(sub_45_carry[14]), .Y(N145) );
  AND2X1 U238 ( .A(n135), .B(n136), .Y(sub_45_carry[14]) );
  XOR2X1 U239 ( .A(n136), .B(n135), .Y(N144) );
endmodule

