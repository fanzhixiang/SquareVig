##
## LEF for PtnCells ;
## created by Encounter v10.13-s272_1 on Thu May 19 19:49:16 2016
##

VERSION 5.6 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO gcd
  CLASS BLOCK ;
  SIZE 97.1700 BY 90.6400 ;
  FOREIGN gcd 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN A_in[7] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT -0.1400 90.5000 0.1400 90.7800 ;
    END
  END A_in[7]
  PIN A_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8888 LAYER METAL3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.0076 LAYER METAL3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.63 LAYER METAL3  ;
    ANTENNAMAXAREACAR 24.8598 LAYER METAL3  ;
    ANTENNAMAXSIDEAREACAR 95.0831 LAYER METAL3  ;
    ANTENNAMAXCUTCAR 0.357672 LAYER VIA34  ;
    PORT
      LAYER METAL3 ;
        RECT 0.0000 77.5500 0.7300 77.8300 ;
    END
  END A_in[6]
  PIN A_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2568 LAYER METAL3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6274 LAYER METAL3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.63 LAYER METAL3  ;
    ANTENNAMAXAREACAR 14.2776 LAYER METAL3  ;
    ANTENNAMAXSIDEAREACAR 55.1263 LAYER METAL3  ;
    ANTENNAMAXCUTCAR 0.500741 LAYER VIA34  ;
    PORT
      LAYER METAL3 ;
        RECT 0.0000 64.6000 0.7300 64.8800 ;
    END
  END A_in[5]
  PIN A_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1183 LAYER METAL3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3715 LAYER METAL3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.63 LAYER METAL3  ;
    ANTENNAMAXAREACAR 13.7367 LAYER METAL3  ;
    ANTENNAMAXSIDEAREACAR 53.3589 LAYER METAL3  ;
    ANTENNAMAXCUTCAR 0.357672 LAYER VIA34  ;
    PORT
      LAYER METAL3 ;
        RECT 0.0000 51.6550 0.7300 51.9350 ;
    END
  END A_in[4]
  PIN A_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8953 LAYER METAL3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.2441 LAYER METAL3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.63 LAYER METAL3  ;
    ANTENNAMAXAREACAR 13.13 LAYER METAL3  ;
    ANTENNAMAXSIDEAREACAR 51.5811 LAYER METAL3  ;
    ANTENNAMAXCUTCAR 0.500741 LAYER VIA34  ;
    PORT
      LAYER METAL3 ;
        RECT 0.0000 38.7050 0.7300 38.9850 ;
    END
  END A_in[3]
  PIN A_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.3522 LAYER METAL3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.7619 LAYER METAL3  ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34  ;
    ANTENNAPARTIALMETALAREA 1.7024 LAYER METAL4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7416 LAYER METAL4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.63 LAYER METAL4  ;
    ANTENNAMAXAREACAR 7.91463 LAYER METAL4  ;
    ANTENNAMAXSIDEAREACAR 32.8965 LAYER METAL4  ;
    ANTENNAMAXCUTCAR 0.608042 LAYER VIA45  ;
    PORT
      LAYER METAL3 ;
        RECT 0.0000 25.7550 0.7300 26.0350 ;
    END
  END A_in[2]
  PIN A_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8266 LAYER METAL3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.494 LAYER METAL3  ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA34  ;
    ANTENNAPARTIALMETALAREA 0.2352 LAYER METAL4  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1872 LAYER METAL4  ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER VIA45  ;
    ANTENNAPARTIALMETALAREA 11.0096 LAYER METAL5  ;
    ANTENNAPARTIALMETALSIDEAREA 41.976 LAYER METAL5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.63 LAYER METAL5  ;
    ANTENNAMAXAREACAR 28.324 LAYER METAL5  ;
    ANTENNAMAXSIDEAREACAR 110.162 LAYER METAL5  ;
    PORT
      LAYER METAL3 ;
        RECT 0.0000 12.8100 0.7300 13.0900 ;
    END
  END A_in[1]
  PIN A_in[0] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT -0.1400 -0.1400 0.1400 0.1400 ;
    END
  END A_in[0]
  PIN B_in[7] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 97.0250 90.5000 97.3050 90.7800 ;
    END
  END B_in[7]
  PIN B_in[6] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 83.1450 90.5000 83.4250 90.7800 ;
    END
  END B_in[6]
  PIN B_in[5] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 69.2650 90.5000 69.5450 90.7800 ;
    END
  END B_in[5]
  PIN B_in[4] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 55.3850 90.5000 55.6650 90.7800 ;
    END
  END B_in[4]
  PIN B_in[3] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 41.5050 90.5000 41.7850 90.7800 ;
    END
  END B_in[3]
  PIN B_in[2] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 27.6200 90.5000 27.9000 90.7800 ;
    END
  END B_in[2]
  PIN B_in[1] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 13.7400 90.5000 14.0200 90.7800 ;
    END
  END B_in[1]
  PIN B_in[0] 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT -0.1400 90.5000 0.1400 90.7800 ;
    END
  END B_in[0]
  PIN clk 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT -0.1400 -0.1400 0.1400 0.1400 ;
    END
  END clk
  PIN rst_n 
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 48.4450 -0.1400 48.7250 0.1400 ;
    END
  END rst_n
  PIN out[7] 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.0300 90.5000 97.3100 90.7800 ;
    END
  END out[7]
  PIN out[6] 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.0300 77.5500 97.3100 77.8300 ;
    END
  END out[6]
  PIN out[5] 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.0300 64.6000 97.3100 64.8800 ;
    END
  END out[5]
  PIN out[4] 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.0300 51.6550 97.3100 51.9350 ;
    END
  END out[4]
  PIN out[3] 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.0300 38.7050 97.3100 38.9850 ;
    END
  END out[3]
  PIN out[2] 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.0300 25.7550 97.3100 26.0350 ;
    END
  END out[2]
  PIN out[1] 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.0300 12.8100 97.3100 13.0900 ;
    END
  END out[1]
  PIN out[0] 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL3 ;
        RECT 97.0300 -0.1400 97.3100 0.1400 ;
    END
  END out[0]
  PIN done 
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL2 ;
        RECT 97.0300 -0.1400 97.3100 0.1400 ;
    END
  END done
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER METAL5 ;
        RECT 0.0000 81.2200 2.0000 83.2200 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 95.1700 81.2200 97.1700 83.2200 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 3.1400 0.0000 5.1400 2.0000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 3.1400 88.6400 5.1400 90.6400 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 92.2850 0.0000 94.2850 2.0000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 92.2850 88.6400 94.2850 90.6400 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 0.0000 2.9000 2.0000 4.9000 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 95.1700 2.9000 97.1700 4.9000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 7.7000 0.0000 9.7000 2.0000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 7.7000 88.6400 9.7000 90.6400 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 87.7250 0.0000 89.7250 2.0000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 87.7250 88.6400 89.7250 90.6400 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 0.0000 7.4600 2.0000 9.4600 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 95.1700 7.4600 97.1700 9.4600 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 0.0000 85.7800 2.0000 87.7800 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 95.1700 85.7800 97.1700 87.7800 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER METAL5 ;
        RECT 0.0000 83.5000 2.0000 85.5000 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 95.1700 83.5000 97.1700 85.5000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 0.8600 0.0000 2.8600 2.0000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 0.8600 88.6400 2.8600 90.6400 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 94.5650 0.0000 96.5650 2.0000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 94.5650 88.6400 96.5650 90.6400 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 0.0000 0.6200 2.0000 2.6200 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 95.1700 0.6200 97.1700 2.6200 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 5.4200 0.0000 7.4200 2.0000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 5.4200 88.6400 7.4200 90.6400 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 90.0050 0.0000 92.0050 2.0000 ;
    END
    PORT
      LAYER METAL4 ;
        RECT 90.0050 88.6400 92.0050 90.6400 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 0.0000 5.1800 2.0000 7.1800 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 95.1700 5.1800 97.1700 7.1800 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 0.0000 88.0600 2.0000 90.0600 ;
    END
    PORT
      LAYER METAL5 ;
        RECT 95.1700 88.0600 97.1700 90.0600 ;
    END
  END VSS
  OBS
    LAYER METAL1 ;
      RECT 0.0000 0.0000 97.1700 90.6400 ;
    LAYER METAL2 ;
      RECT 0.0000 0.0000 97.1700 90.6400 ;
    LAYER METAL3 ;
      RECT 0.4200 90.2200 97.1700 90.6400 ;
      RECT 0.0000 78.1100 97.1700 90.2200 ;
      RECT 1.0100 77.2700 97.1700 78.1100 ;
      RECT 0.0000 65.1600 97.1700 77.2700 ;
      RECT 1.0100 64.3200 97.1700 65.1600 ;
      RECT 0.0000 52.2150 97.1700 64.3200 ;
      RECT 1.0100 51.3750 97.1700 52.2150 ;
      RECT 0.0000 39.2650 97.1700 51.3750 ;
      RECT 1.0100 38.4250 97.1700 39.2650 ;
      RECT 0.0000 26.3150 97.1700 38.4250 ;
      RECT 1.0100 25.4750 97.1700 26.3150 ;
      RECT 0.0000 0.0000 97.1700 25.4750 ;
